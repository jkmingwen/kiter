library ieee;
use ieee.std_logic_1164.all;

$ENTITY_DECLARATION

-- architecture Behavioral of const_value_$N_OUTPUTS is
architecture Behavioral of $COMPONENT_NAME is
begin

$PROCESS_BEHAVIOUR

end Behavioral;
