-- Broadcast
-- Takes in 1 input data and sends to all output ports

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

$ENTITY_DECLARATION

architecture Behavioral of $COMPONENT_NAME is

begin

    $PROCESS_BEHAVIOUR

end Behavioral;
