--------------------------------------------------------------------------------
--                         Compressor_6_3_F125_uid69
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_F125_uid69 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_F125_uid69 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <=
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         Compressor_14_3_F125_uid79
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_F125_uid79 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_F125_uid79 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <=
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        Compressor_23_3_F125_uid193
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_F125_uid193 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_F125_uid193 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <=
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         Compressor_3_2_F125_uid223
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_F125_uid223 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_F125_uid223 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <=
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x19_F125_uid6
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x19_F125_uid6 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(18 downto 0);
          R : out  std_logic_vector(35 downto 0)   );
end entity;

architecture arch of DSPBlock_17x19_F125_uid6 is
signal Mint :  std_logic_vector(35 downto 0);
signal M :  std_logic_vector(35 downto 0);
signal Rtmp :  std_logic_vector(35 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(35 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_19x1_F125_uid8
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_19x1_F125_uid8 is
    port (clk : in std_logic;
          X : in  std_logic_vector(18 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(18 downto 0)   );
end entity;

architecture arch of DSPBlock_19x1_F125_uid8 is
signal Mint :  std_logic_vector(19 downto 0);
signal M :  std_logic_vector(18 downto 0);
signal Rtmp :  std_logic_vector(18 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(18 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_18x1_F125_uid10
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_18x1_F125_uid10 is
    port (clk : in std_logic;
          X : in  std_logic_vector(17 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(17 downto 0)   );
end entity;

architecture arch of DSPBlock_18x1_F125_uid10 is
signal Mint :  std_logic_vector(18 downto 0);
signal M :  std_logic_vector(17 downto 0);
signal Rtmp :  std_logic_vector(17 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(17 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x18_F125_uid12
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x18_F125_uid12 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(17 downto 0);
          R : out  std_logic_vector(17 downto 0)   );
end entity;

architecture arch of DSPBlock_1x18_F125_uid12 is
signal Mint :  std_logic_vector(18 downto 0);
signal M :  std_logic_vector(17 downto 0);
signal Rtmp :  std_logic_vector(17 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(17 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x17_F125_uid14
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x17_F125_uid14 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(16 downto 0);
          R : out  std_logic_vector(16 downto 0)   );
end entity;

architecture arch of DSPBlock_1x17_F125_uid14 is
signal Mint :  std_logic_vector(17 downto 0);
signal M :  std_logic_vector(16 downto 0);
signal Rtmp :  std_logic_vector(16 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(16 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x1_F125_uid16
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x1_F125_uid16 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(16 downto 0)   );
end entity;

architecture arch of DSPBlock_17x1_F125_uid16 is
signal Mint :  std_logic_vector(17 downto 0);
signal M :  std_logic_vector(16 downto 0);
signal Rtmp :  std_logic_vector(16 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(16 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_16x1_F125_uid18
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_16x1_F125_uid18 is
    port (clk : in std_logic;
          X : in  std_logic_vector(15 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(15 downto 0)   );
end entity;

architecture arch of DSPBlock_16x1_F125_uid18 is
signal Mint :  std_logic_vector(16 downto 0);
signal M :  std_logic_vector(15 downto 0);
signal Rtmp :  std_logic_vector(15 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(15 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x16_F125_uid20
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x16_F125_uid20 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(15 downto 0);
          R : out  std_logic_vector(15 downto 0)   );
end entity;

architecture arch of DSPBlock_1x16_F125_uid20 is
signal Mint :  std_logic_vector(16 downto 0);
signal M :  std_logic_vector(15 downto 0);
signal Rtmp :  std_logic_vector(15 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(15 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x15_F125_uid22
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x15_F125_uid22 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(14 downto 0);
          R : out  std_logic_vector(14 downto 0)   );
end entity;

architecture arch of DSPBlock_1x15_F125_uid22 is
signal Mint :  std_logic_vector(15 downto 0);
signal M :  std_logic_vector(14 downto 0);
signal Rtmp :  std_logic_vector(14 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(14 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_15x1_F125_uid24
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_15x1_F125_uid24 is
    port (clk : in std_logic;
          X : in  std_logic_vector(14 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(14 downto 0)   );
end entity;

architecture arch of DSPBlock_15x1_F125_uid24 is
signal Mint :  std_logic_vector(15 downto 0);
signal M :  std_logic_vector(14 downto 0);
signal Rtmp :  std_logic_vector(14 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(14 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_14x1_F125_uid26
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_14x1_F125_uid26 is
    port (clk : in std_logic;
          X : in  std_logic_vector(13 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(13 downto 0)   );
end entity;

architecture arch of DSPBlock_14x1_F125_uid26 is
signal Mint :  std_logic_vector(14 downto 0);
signal M :  std_logic_vector(13 downto 0);
signal Rtmp :  std_logic_vector(13 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(13 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x14_F125_uid28
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x14_F125_uid28 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(13 downto 0);
          R : out  std_logic_vector(13 downto 0)   );
end entity;

architecture arch of DSPBlock_1x14_F125_uid28 is
signal Mint :  std_logic_vector(14 downto 0);
signal M :  std_logic_vector(13 downto 0);
signal Rtmp :  std_logic_vector(13 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(13 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_13x1_F125_uid30
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_13x1_F125_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(12 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(12 downto 0)   );
end entity;

architecture arch of DSPBlock_13x1_F125_uid30 is
signal Mint :  std_logic_vector(13 downto 0);
signal M :  std_logic_vector(12 downto 0);
signal Rtmp :  std_logic_vector(12 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(12 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x13_F125_uid32
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x13_F125_uid32 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(12 downto 0);
          R : out  std_logic_vector(12 downto 0)   );
end entity;

architecture arch of DSPBlock_1x13_F125_uid32 is
signal Mint :  std_logic_vector(13 downto 0);
signal M :  std_logic_vector(12 downto 0);
signal Rtmp :  std_logic_vector(12 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(12 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x12_F125_uid34
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x12_F125_uid34 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(11 downto 0);
          R : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of DSPBlock_1x12_F125_uid34 is
signal Mint :  std_logic_vector(12 downto 0);
signal M :  std_logic_vector(11 downto 0);
signal Rtmp :  std_logic_vector(11 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(11 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_12x1_F125_uid36
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_12x1_F125_uid36 is
    port (clk : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of DSPBlock_12x1_F125_uid36 is
signal Mint :  std_logic_vector(12 downto 0);
signal M :  std_logic_vector(11 downto 0);
signal Rtmp :  std_logic_vector(11 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(11 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_11x1_F125_uid38
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_11x1_F125_uid38 is
    port (clk : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(10 downto 0)   );
end entity;

architecture arch of DSPBlock_11x1_F125_uid38 is
signal Mint :  std_logic_vector(11 downto 0);
signal M :  std_logic_vector(10 downto 0);
signal Rtmp :  std_logic_vector(10 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(10 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x11_F125_uid40
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x11_F125_uid40 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(10 downto 0);
          R : out  std_logic_vector(10 downto 0)   );
end entity;

architecture arch of DSPBlock_1x11_F125_uid40 is
signal Mint :  std_logic_vector(11 downto 0);
signal M :  std_logic_vector(10 downto 0);
signal Rtmp :  std_logic_vector(10 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(10 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_10x1_F125_uid42
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_10x1_F125_uid42 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of DSPBlock_10x1_F125_uid42 is
signal Mint :  std_logic_vector(10 downto 0);
signal M :  std_logic_vector(9 downto 0);
signal Rtmp :  std_logic_vector(9 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(9 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x10_F125_uid44
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x10_F125_uid44 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(9 downto 0);
          R : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of DSPBlock_1x10_F125_uid44 is
signal Mint :  std_logic_vector(10 downto 0);
signal M :  std_logic_vector(9 downto 0);
signal Rtmp :  std_logic_vector(9 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(9 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_9x1_F125_uid46
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_9x1_F125_uid46 is
    port (clk : in std_logic;
          X : in  std_logic_vector(8 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of DSPBlock_9x1_F125_uid46 is
signal Mint :  std_logic_vector(9 downto 0);
signal M :  std_logic_vector(8 downto 0);
signal Rtmp :  std_logic_vector(8 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(8 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x9_F125_uid48
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x9_F125_uid48 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(8 downto 0);
          R : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of DSPBlock_1x9_F125_uid48 is
signal Mint :  std_logic_vector(9 downto 0);
signal M :  std_logic_vector(8 downto 0);
signal Rtmp :  std_logic_vector(8 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(8 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_8x1_F125_uid50
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_8x1_F125_uid50 is
    port (clk : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(7 downto 0)   );
end entity;

architecture arch of DSPBlock_8x1_F125_uid50 is
signal Mint :  std_logic_vector(8 downto 0);
signal M :  std_logic_vector(7 downto 0);
signal Rtmp :  std_logic_vector(7 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(7 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x8_F125_uid52
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x8_F125_uid52 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(7 downto 0)   );
end entity;

architecture arch of DSPBlock_1x8_F125_uid52 is
signal Mint :  std_logic_vector(8 downto 0);
signal M :  std_logic_vector(7 downto 0);
signal Rtmp :  std_logic_vector(7 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(7 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_7x1_F125_uid54
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_7x1_F125_uid54 is
    port (clk : in std_logic;
          X : in  std_logic_vector(6 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of DSPBlock_7x1_F125_uid54 is
signal Mint :  std_logic_vector(7 downto 0);
signal M :  std_logic_vector(6 downto 0);
signal Rtmp :  std_logic_vector(6 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(6 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x7_F125_uid56
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x7_F125_uid56 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(6 downto 0);
          R : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of DSPBlock_1x7_F125_uid56 is
signal Mint :  std_logic_vector(7 downto 0);
signal M :  std_logic_vector(6 downto 0);
signal Rtmp :  std_logic_vector(6 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(6 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x6_F125_uid58
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x6_F125_uid58 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of DSPBlock_1x6_F125_uid58 is
signal Mint :  std_logic_vector(6 downto 0);
signal M :  std_logic_vector(5 downto 0);
signal Rtmp :  std_logic_vector(5 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(5 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_1x5_F125_uid60
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_1x5_F125_uid60 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of DSPBlock_1x5_F125_uid60 is
signal Mint :  std_logic_vector(5 downto 0);
signal M :  std_logic_vector(4 downto 0);
signal Rtmp :  std_logic_vector(4 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(4 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_5x1_F125_uid62
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_5x1_F125_uid62 is
    port (clk : in std_logic;
          X : in  std_logic_vector(4 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of DSPBlock_5x1_F125_uid62 is
signal Mint :  std_logic_vector(5 downto 0);
signal M :  std_logic_vector(4 downto 0);
signal Rtmp :  std_logic_vector(4 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(4 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_4x1_F125_uid64
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_4x1_F125_uid64 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of DSPBlock_4x1_F125_uid64 is
signal Mint :  std_logic_vector(4 downto 0);
signal M :  std_logic_vector(3 downto 0);
signal Rtmp :  std_logic_vector(3 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(3 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_3x19_F125_uid66
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors:
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_3x19_F125_uid66 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(18 downto 0);
          R : out  std_logic_vector(21 downto 0)   );
end entity;

architecture arch of DSPBlock_3x19_F125_uid66 is
signal Mint :  std_logic_vector(21 downto 0);
signal M :  std_logic_vector(21 downto 0);
signal Rtmp :  std_logic_vector(21 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(21 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_64_F125_uid443
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_64_F125_uid443 is
    port (clk : in std_logic;
          X : in  std_logic_vector(63 downto 0);
          Y : in  std_logic_vector(63 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(63 downto 0)   );
end entity;

architecture arch of IntAdder_64_F125_uid443 is
signal Rtmp :  std_logic_vector(63 downto 0);
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          IntMultiplier_F125_uid2
-- VHDL generated for Zynq7000 @ 125MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 8
-- Target frequency (MHz): 125
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_F125_uid2 is
    port (clk : in std_logic;
          X : in  std_logic_vector(33 downto 0);
          Y : in  std_logic_vector(33 downto 0);
          R : out  std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntMultiplier_F125_uid2 is
   component DSPBlock_17x19_F125_uid6 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(18 downto 0);
             R : out  std_logic_vector(35 downto 0)   );
   end component;

   component DSPBlock_19x1_F125_uid8 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(18 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(18 downto 0)   );
   end component;

   component DSPBlock_18x1_F125_uid10 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(17 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(17 downto 0)   );
   end component;

   component DSPBlock_1x18_F125_uid12 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(17 downto 0);
             R : out  std_logic_vector(17 downto 0)   );
   end component;

   component DSPBlock_1x17_F125_uid14 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(16 downto 0);
             R : out  std_logic_vector(16 downto 0)   );
   end component;

   component DSPBlock_17x1_F125_uid16 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(16 downto 0)   );
   end component;

   component DSPBlock_16x1_F125_uid18 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(15 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(15 downto 0)   );
   end component;

   component DSPBlock_1x16_F125_uid20 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(15 downto 0);
             R : out  std_logic_vector(15 downto 0)   );
   end component;

   component DSPBlock_1x15_F125_uid22 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(14 downto 0);
             R : out  std_logic_vector(14 downto 0)   );
   end component;

   component DSPBlock_15x1_F125_uid24 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(14 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(14 downto 0)   );
   end component;

   component DSPBlock_14x1_F125_uid26 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(13 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(13 downto 0)   );
   end component;

   component DSPBlock_1x14_F125_uid28 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(13 downto 0);
             R : out  std_logic_vector(13 downto 0)   );
   end component;

   component DSPBlock_13x1_F125_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(12 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(12 downto 0)   );
   end component;

   component DSPBlock_1x13_F125_uid32 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(12 downto 0);
             R : out  std_logic_vector(12 downto 0)   );
   end component;

   component DSPBlock_1x12_F125_uid34 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(11 downto 0);
             R : out  std_logic_vector(11 downto 0)   );
   end component;

   component DSPBlock_12x1_F125_uid36 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(11 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(11 downto 0)   );
   end component;

   component DSPBlock_11x1_F125_uid38 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(10 downto 0)   );
   end component;

   component DSPBlock_1x11_F125_uid40 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(10 downto 0);
             R : out  std_logic_vector(10 downto 0)   );
   end component;

   component DSPBlock_10x1_F125_uid42 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(9 downto 0)   );
   end component;

   component DSPBlock_1x10_F125_uid44 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(9 downto 0);
             R : out  std_logic_vector(9 downto 0)   );
   end component;

   component DSPBlock_9x1_F125_uid46 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(8 downto 0)   );
   end component;

   component DSPBlock_1x9_F125_uid48 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(8 downto 0);
             R : out  std_logic_vector(8 downto 0)   );
   end component;

   component DSPBlock_8x1_F125_uid50 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(7 downto 0)   );
   end component;

   component DSPBlock_1x8_F125_uid52 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(7 downto 0)   );
   end component;

   component DSPBlock_7x1_F125_uid54 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(6 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(6 downto 0)   );
   end component;

   component DSPBlock_1x7_F125_uid56 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(6 downto 0);
             R : out  std_logic_vector(6 downto 0)   );
   end component;

   component DSPBlock_1x6_F125_uid58 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(5 downto 0)   );
   end component;

   component DSPBlock_1x5_F125_uid60 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component DSPBlock_5x1_F125_uid62 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(4 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component DSPBlock_4x1_F125_uid64 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component DSPBlock_3x19_F125_uid66 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(18 downto 0);
             R : out  std_logic_vector(21 downto 0)   );
   end component;

   component Compressor_6_3_F125_uid69 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_F125_uid79 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_23_3_F125_uid193 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_F125_uid223 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntAdder_64_F125_uid443 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(63 downto 0);
             Y : in  std_logic_vector(63 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(63 downto 0)   );
   end component;

signal XX_m3 :  std_logic_vector(33 downto 0);
signal YY_m3 :  std_logic_vector(33 downto 0);
signal tile_0_X :  std_logic_vector(16 downto 0);
signal tile_0_Y :  std_logic_vector(18 downto 0);
signal tile_0_output :  std_logic_vector(35 downto 0);
signal tile_0_filtered_output :  unsigned(35-0 downto 0);
signal bh4_w0_0 :  std_logic;
signal bh4_w1_0 :  std_logic;
signal bh4_w2_0 :  std_logic;
signal bh4_w3_0 :  std_logic;
signal bh4_w4_0 :  std_logic;
signal bh4_w5_0 :  std_logic;
signal bh4_w6_0 :  std_logic;
signal bh4_w7_0 :  std_logic;
signal bh4_w8_0 :  std_logic;
signal bh4_w9_0 :  std_logic;
signal bh4_w10_0 :  std_logic;
signal bh4_w11_0 :  std_logic;
signal bh4_w12_0 :  std_logic;
signal bh4_w13_0 :  std_logic;
signal bh4_w14_0 :  std_logic;
signal bh4_w15_0 :  std_logic;
signal bh4_w16_0 :  std_logic;
signal bh4_w17_0 :  std_logic;
signal bh4_w18_0 :  std_logic;
signal bh4_w19_0 :  std_logic;
signal bh4_w20_0 :  std_logic;
signal bh4_w21_0 :  std_logic;
signal bh4_w22_0 :  std_logic;
signal bh4_w23_0 :  std_logic;
signal bh4_w24_0 :  std_logic;
signal bh4_w25_0 :  std_logic;
signal bh4_w26_0 :  std_logic;
signal bh4_w27_0 :  std_logic;
signal bh4_w28_0 :  std_logic;
signal bh4_w29_0 :  std_logic;
signal bh4_w30_0 :  std_logic;
signal bh4_w31_0 :  std_logic;
signal bh4_w32_0 :  std_logic;
signal bh4_w33_0 :  std_logic;
signal bh4_w34_0 :  std_logic;
signal bh4_w35_0 :  std_logic;
signal tile_1_X :  std_logic_vector(18 downto 0);
signal tile_1_Y :  std_logic_vector(0 downto 0);
signal tile_1_output :  std_logic_vector(18 downto 0);
signal tile_1_filtered_output :  unsigned(18-0 downto 0);
signal bh4_w0_1 :  std_logic;
signal bh4_w1_1 :  std_logic;
signal bh4_w2_1 :  std_logic;
signal bh4_w3_1 :  std_logic;
signal bh4_w4_1 :  std_logic;
signal bh4_w5_1 :  std_logic;
signal bh4_w6_1 :  std_logic;
signal bh4_w7_1 :  std_logic;
signal bh4_w8_1 :  std_logic;
signal bh4_w9_1 :  std_logic;
signal bh4_w10_1 :  std_logic;
signal bh4_w11_1 :  std_logic;
signal bh4_w12_1 :  std_logic;
signal bh4_w13_1 :  std_logic;
signal bh4_w14_1 :  std_logic;
signal bh4_w15_1 :  std_logic;
signal bh4_w16_1 :  std_logic;
signal bh4_w17_1 :  std_logic;
signal bh4_w18_1 :  std_logic;
signal tile_2_X :  std_logic_vector(17 downto 0);
signal tile_2_Y :  std_logic_vector(0 downto 0);
signal tile_2_output :  std_logic_vector(17 downto 0);
signal tile_2_filtered_output :  unsigned(17-0 downto 0);
signal bh4_w0_2 :  std_logic;
signal bh4_w1_2 :  std_logic;
signal bh4_w2_2 :  std_logic;
signal bh4_w3_2 :  std_logic;
signal bh4_w4_2 :  std_logic;
signal bh4_w5_2 :  std_logic;
signal bh4_w6_2 :  std_logic;
signal bh4_w7_2 :  std_logic;
signal bh4_w8_2 :  std_logic;
signal bh4_w9_2 :  std_logic;
signal bh4_w10_2 :  std_logic;
signal bh4_w11_2 :  std_logic;
signal bh4_w12_2 :  std_logic;
signal bh4_w13_2 :  std_logic;
signal bh4_w14_2 :  std_logic;
signal bh4_w15_2 :  std_logic;
signal bh4_w16_2 :  std_logic;
signal bh4_w17_2 :  std_logic;
signal tile_3_X :  std_logic_vector(0 downto 0);
signal tile_3_Y :  std_logic_vector(17 downto 0);
signal tile_3_output :  std_logic_vector(17 downto 0);
signal tile_3_filtered_output :  unsigned(17-0 downto 0);
signal bh4_w0_3 :  std_logic;
signal bh4_w1_3 :  std_logic;
signal bh4_w2_3 :  std_logic;
signal bh4_w3_3 :  std_logic;
signal bh4_w4_3 :  std_logic;
signal bh4_w5_3 :  std_logic;
signal bh4_w6_3 :  std_logic;
signal bh4_w7_3 :  std_logic;
signal bh4_w8_3 :  std_logic;
signal bh4_w9_3 :  std_logic;
signal bh4_w10_3 :  std_logic;
signal bh4_w11_3 :  std_logic;
signal bh4_w12_3 :  std_logic;
signal bh4_w13_3 :  std_logic;
signal bh4_w14_3 :  std_logic;
signal bh4_w15_3 :  std_logic;
signal bh4_w16_3 :  std_logic;
signal bh4_w17_3 :  std_logic;
signal tile_4_X :  std_logic_vector(0 downto 0);
signal tile_4_Y :  std_logic_vector(16 downto 0);
signal tile_4_output :  std_logic_vector(16 downto 0);
signal tile_4_filtered_output :  unsigned(16-0 downto 0);
signal bh4_w0_4 :  std_logic;
signal bh4_w1_4 :  std_logic;
signal bh4_w2_4 :  std_logic;
signal bh4_w3_4 :  std_logic;
signal bh4_w4_4 :  std_logic;
signal bh4_w5_4 :  std_logic;
signal bh4_w6_4 :  std_logic;
signal bh4_w7_4 :  std_logic;
signal bh4_w8_4 :  std_logic;
signal bh4_w9_4 :  std_logic;
signal bh4_w10_4 :  std_logic;
signal bh4_w11_4 :  std_logic;
signal bh4_w12_4 :  std_logic;
signal bh4_w13_4 :  std_logic;
signal bh4_w14_4 :  std_logic;
signal bh4_w15_4 :  std_logic;
signal bh4_w16_4 :  std_logic;
signal tile_5_X :  std_logic_vector(16 downto 0);
signal tile_5_Y :  std_logic_vector(0 downto 0);
signal tile_5_output :  std_logic_vector(16 downto 0);
signal tile_5_filtered_output :  unsigned(16-0 downto 0);
signal bh4_w0_5 :  std_logic;
signal bh4_w1_5 :  std_logic;
signal bh4_w2_5 :  std_logic;
signal bh4_w3_5 :  std_logic;
signal bh4_w4_5 :  std_logic;
signal bh4_w5_5 :  std_logic;
signal bh4_w6_5 :  std_logic;
signal bh4_w7_5 :  std_logic;
signal bh4_w8_5 :  std_logic;
signal bh4_w9_5 :  std_logic;
signal bh4_w10_5 :  std_logic;
signal bh4_w11_5 :  std_logic;
signal bh4_w12_5 :  std_logic;
signal bh4_w13_5 :  std_logic;
signal bh4_w14_5 :  std_logic;
signal bh4_w15_5 :  std_logic;
signal bh4_w16_5 :  std_logic;
signal tile_6_X :  std_logic_vector(15 downto 0);
signal tile_6_Y :  std_logic_vector(0 downto 0);
signal tile_6_output :  std_logic_vector(15 downto 0);
signal tile_6_filtered_output :  unsigned(15-0 downto 0);
signal bh4_w0_6 :  std_logic;
signal bh4_w1_6 :  std_logic;
signal bh4_w2_6 :  std_logic;
signal bh4_w3_6 :  std_logic;
signal bh4_w4_6 :  std_logic;
signal bh4_w5_6 :  std_logic;
signal bh4_w6_6 :  std_logic;
signal bh4_w7_6 :  std_logic;
signal bh4_w8_6 :  std_logic;
signal bh4_w9_6 :  std_logic;
signal bh4_w10_6 :  std_logic;
signal bh4_w11_6 :  std_logic;
signal bh4_w12_6 :  std_logic;
signal bh4_w13_6 :  std_logic;
signal bh4_w14_6 :  std_logic;
signal bh4_w15_6 :  std_logic;
signal tile_7_X :  std_logic_vector(0 downto 0);
signal tile_7_Y :  std_logic_vector(15 downto 0);
signal tile_7_output :  std_logic_vector(15 downto 0);
signal tile_7_filtered_output :  unsigned(15-0 downto 0);
signal bh4_w0_7 :  std_logic;
signal bh4_w1_7 :  std_logic;
signal bh4_w2_7 :  std_logic;
signal bh4_w3_7 :  std_logic;
signal bh4_w4_7 :  std_logic;
signal bh4_w5_7 :  std_logic;
signal bh4_w6_7 :  std_logic;
signal bh4_w7_7 :  std_logic;
signal bh4_w8_7 :  std_logic;
signal bh4_w9_7 :  std_logic;
signal bh4_w10_7 :  std_logic;
signal bh4_w11_7 :  std_logic;
signal bh4_w12_7 :  std_logic;
signal bh4_w13_7 :  std_logic;
signal bh4_w14_7 :  std_logic;
signal bh4_w15_7 :  std_logic;
signal tile_8_X :  std_logic_vector(0 downto 0);
signal tile_8_Y :  std_logic_vector(14 downto 0);
signal tile_8_output :  std_logic_vector(14 downto 0);
signal tile_8_filtered_output :  unsigned(14-0 downto 0);
signal bh4_w0_8 :  std_logic;
signal bh4_w1_8 :  std_logic;
signal bh4_w2_8 :  std_logic;
signal bh4_w3_8 :  std_logic;
signal bh4_w4_8 :  std_logic;
signal bh4_w5_8 :  std_logic;
signal bh4_w6_8 :  std_logic;
signal bh4_w7_8 :  std_logic;
signal bh4_w8_8 :  std_logic;
signal bh4_w9_8 :  std_logic;
signal bh4_w10_8 :  std_logic;
signal bh4_w11_8 :  std_logic;
signal bh4_w12_8 :  std_logic;
signal bh4_w13_8 :  std_logic;
signal bh4_w14_8 :  std_logic;
signal tile_9_X :  std_logic_vector(14 downto 0);
signal tile_9_Y :  std_logic_vector(0 downto 0);
signal tile_9_output :  std_logic_vector(14 downto 0);
signal tile_9_filtered_output :  unsigned(14-0 downto 0);
signal bh4_w0_9 :  std_logic;
signal bh4_w1_9 :  std_logic;
signal bh4_w2_9 :  std_logic;
signal bh4_w3_9 :  std_logic;
signal bh4_w4_9 :  std_logic;
signal bh4_w5_9 :  std_logic;
signal bh4_w6_9 :  std_logic;
signal bh4_w7_9 :  std_logic;
signal bh4_w8_9 :  std_logic;
signal bh4_w9_9 :  std_logic;
signal bh4_w10_9 :  std_logic;
signal bh4_w11_9 :  std_logic;
signal bh4_w12_9 :  std_logic;
signal bh4_w13_9 :  std_logic;
signal bh4_w14_9 :  std_logic;
signal tile_10_X :  std_logic_vector(13 downto 0);
signal tile_10_Y :  std_logic_vector(0 downto 0);
signal tile_10_output :  std_logic_vector(13 downto 0);
signal tile_10_filtered_output :  unsigned(13-0 downto 0);
signal bh4_w0_10 :  std_logic;
signal bh4_w1_10 :  std_logic;
signal bh4_w2_10 :  std_logic;
signal bh4_w3_10 :  std_logic;
signal bh4_w4_10 :  std_logic;
signal bh4_w5_10 :  std_logic;
signal bh4_w6_10 :  std_logic;
signal bh4_w7_10 :  std_logic;
signal bh4_w8_10 :  std_logic;
signal bh4_w9_10 :  std_logic;
signal bh4_w10_10 :  std_logic;
signal bh4_w11_10 :  std_logic;
signal bh4_w12_10 :  std_logic;
signal bh4_w13_10 :  std_logic;
signal tile_11_X :  std_logic_vector(0 downto 0);
signal tile_11_Y :  std_logic_vector(13 downto 0);
signal tile_11_output :  std_logic_vector(13 downto 0);
signal tile_11_filtered_output :  unsigned(13-0 downto 0);
signal bh4_w0_11 :  std_logic;
signal bh4_w1_11 :  std_logic;
signal bh4_w2_11 :  std_logic;
signal bh4_w3_11 :  std_logic;
signal bh4_w4_11 :  std_logic;
signal bh4_w5_11 :  std_logic;
signal bh4_w6_11 :  std_logic;
signal bh4_w7_11 :  std_logic;
signal bh4_w8_11 :  std_logic;
signal bh4_w9_11 :  std_logic;
signal bh4_w10_11 :  std_logic;
signal bh4_w11_11 :  std_logic;
signal bh4_w12_11 :  std_logic;
signal bh4_w13_11 :  std_logic;
signal tile_12_X :  std_logic_vector(12 downto 0);
signal tile_12_Y :  std_logic_vector(0 downto 0);
signal tile_12_output :  std_logic_vector(12 downto 0);
signal tile_12_filtered_output :  unsigned(12-0 downto 0);
signal bh4_w0_12 :  std_logic;
signal bh4_w1_12 :  std_logic;
signal bh4_w2_12 :  std_logic;
signal bh4_w3_12 :  std_logic;
signal bh4_w4_12 :  std_logic;
signal bh4_w5_12 :  std_logic;
signal bh4_w6_12 :  std_logic;
signal bh4_w7_12 :  std_logic;
signal bh4_w8_12 :  std_logic;
signal bh4_w9_12 :  std_logic;
signal bh4_w10_12 :  std_logic;
signal bh4_w11_12 :  std_logic;
signal bh4_w12_12 :  std_logic;
signal tile_13_X :  std_logic_vector(0 downto 0);
signal tile_13_Y :  std_logic_vector(12 downto 0);
signal tile_13_output :  std_logic_vector(12 downto 0);
signal tile_13_filtered_output :  unsigned(12-0 downto 0);
signal bh4_w0_13 :  std_logic;
signal bh4_w1_13 :  std_logic;
signal bh4_w2_13 :  std_logic;
signal bh4_w3_13 :  std_logic;
signal bh4_w4_13 :  std_logic;
signal bh4_w5_13 :  std_logic;
signal bh4_w6_13 :  std_logic;
signal bh4_w7_13 :  std_logic;
signal bh4_w8_13 :  std_logic;
signal bh4_w9_13 :  std_logic;
signal bh4_w10_13 :  std_logic;
signal bh4_w11_13 :  std_logic;
signal bh4_w12_13 :  std_logic;
signal tile_14_X :  std_logic_vector(0 downto 0);
signal tile_14_Y :  std_logic_vector(11 downto 0);
signal tile_14_output :  std_logic_vector(11 downto 0);
signal tile_14_filtered_output :  unsigned(11-0 downto 0);
signal bh4_w0_14 :  std_logic;
signal bh4_w1_14 :  std_logic;
signal bh4_w2_14 :  std_logic;
signal bh4_w3_14 :  std_logic;
signal bh4_w4_14 :  std_logic;
signal bh4_w5_14 :  std_logic;
signal bh4_w6_14 :  std_logic;
signal bh4_w7_14 :  std_logic;
signal bh4_w8_14 :  std_logic;
signal bh4_w9_14 :  std_logic;
signal bh4_w10_14 :  std_logic;
signal bh4_w11_14 :  std_logic;
signal tile_15_X :  std_logic_vector(11 downto 0);
signal tile_15_Y :  std_logic_vector(0 downto 0);
signal tile_15_output :  std_logic_vector(11 downto 0);
signal tile_15_filtered_output :  unsigned(11-0 downto 0);
signal bh4_w0_15 :  std_logic;
signal bh4_w1_15 :  std_logic;
signal bh4_w2_15 :  std_logic;
signal bh4_w3_15 :  std_logic;
signal bh4_w4_15 :  std_logic;
signal bh4_w5_15 :  std_logic;
signal bh4_w6_15 :  std_logic;
signal bh4_w7_15 :  std_logic;
signal bh4_w8_15 :  std_logic;
signal bh4_w9_15 :  std_logic;
signal bh4_w10_15 :  std_logic;
signal bh4_w11_15 :  std_logic;
signal tile_16_X :  std_logic_vector(10 downto 0);
signal tile_16_Y :  std_logic_vector(0 downto 0);
signal tile_16_output :  std_logic_vector(10 downto 0);
signal tile_16_filtered_output :  unsigned(10-0 downto 0);
signal bh4_w0_16 :  std_logic;
signal bh4_w1_16 :  std_logic;
signal bh4_w2_16 :  std_logic;
signal bh4_w3_16 :  std_logic;
signal bh4_w4_16 :  std_logic;
signal bh4_w5_16 :  std_logic;
signal bh4_w6_16 :  std_logic;
signal bh4_w7_16 :  std_logic;
signal bh4_w8_16 :  std_logic;
signal bh4_w9_16 :  std_logic;
signal bh4_w10_16 :  std_logic;
signal tile_17_X :  std_logic_vector(0 downto 0);
signal tile_17_Y :  std_logic_vector(10 downto 0);
signal tile_17_output :  std_logic_vector(10 downto 0);
signal tile_17_filtered_output :  unsigned(10-0 downto 0);
signal bh4_w0_17 :  std_logic;
signal bh4_w1_17 :  std_logic;
signal bh4_w2_17 :  std_logic;
signal bh4_w3_17 :  std_logic;
signal bh4_w4_17 :  std_logic;
signal bh4_w5_17 :  std_logic;
signal bh4_w6_17 :  std_logic;
signal bh4_w7_17 :  std_logic;
signal bh4_w8_17 :  std_logic;
signal bh4_w9_17 :  std_logic;
signal bh4_w10_17 :  std_logic;
signal tile_18_X :  std_logic_vector(9 downto 0);
signal tile_18_Y :  std_logic_vector(0 downto 0);
signal tile_18_output :  std_logic_vector(9 downto 0);
signal tile_18_filtered_output :  unsigned(9-0 downto 0);
signal bh4_w0_18 :  std_logic;
signal bh4_w1_18 :  std_logic;
signal bh4_w2_18 :  std_logic;
signal bh4_w3_18 :  std_logic;
signal bh4_w4_18 :  std_logic;
signal bh4_w5_18 :  std_logic;
signal bh4_w6_18 :  std_logic;
signal bh4_w7_18 :  std_logic;
signal bh4_w8_18 :  std_logic;
signal bh4_w9_18 :  std_logic;
signal tile_19_X :  std_logic_vector(0 downto 0);
signal tile_19_Y :  std_logic_vector(9 downto 0);
signal tile_19_output :  std_logic_vector(9 downto 0);
signal tile_19_filtered_output :  unsigned(9-0 downto 0);
signal bh4_w0_19 :  std_logic;
signal bh4_w1_19 :  std_logic;
signal bh4_w2_19 :  std_logic;
signal bh4_w3_19 :  std_logic;
signal bh4_w4_19 :  std_logic;
signal bh4_w5_19 :  std_logic;
signal bh4_w6_19 :  std_logic;
signal bh4_w7_19 :  std_logic;
signal bh4_w8_19 :  std_logic;
signal bh4_w9_19 :  std_logic;
signal tile_20_X :  std_logic_vector(8 downto 0);
signal tile_20_Y :  std_logic_vector(0 downto 0);
signal tile_20_output :  std_logic_vector(8 downto 0);
signal tile_20_filtered_output :  unsigned(8-0 downto 0);
signal bh4_w0_20 :  std_logic;
signal bh4_w1_20 :  std_logic;
signal bh4_w2_20 :  std_logic;
signal bh4_w3_20 :  std_logic;
signal bh4_w4_20 :  std_logic;
signal bh4_w5_20 :  std_logic;
signal bh4_w6_20 :  std_logic;
signal bh4_w7_20 :  std_logic;
signal bh4_w8_20 :  std_logic;
signal tile_21_X :  std_logic_vector(0 downto 0);
signal tile_21_Y :  std_logic_vector(8 downto 0);
signal tile_21_output :  std_logic_vector(8 downto 0);
signal tile_21_filtered_output :  unsigned(8-0 downto 0);
signal bh4_w0_21 :  std_logic;
signal bh4_w1_21 :  std_logic;
signal bh4_w2_21 :  std_logic;
signal bh4_w3_21 :  std_logic;
signal bh4_w4_21 :  std_logic;
signal bh4_w5_21 :  std_logic;
signal bh4_w6_21 :  std_logic;
signal bh4_w7_21 :  std_logic;
signal bh4_w8_21 :  std_logic;
signal tile_22_X :  std_logic_vector(7 downto 0);
signal tile_22_Y :  std_logic_vector(0 downto 0);
signal tile_22_output :  std_logic_vector(7 downto 0);
signal tile_22_filtered_output :  unsigned(7-0 downto 0);
signal bh4_w0_22 :  std_logic;
signal bh4_w1_22 :  std_logic;
signal bh4_w2_22 :  std_logic;
signal bh4_w3_22 :  std_logic;
signal bh4_w4_22 :  std_logic;
signal bh4_w5_22 :  std_logic;
signal bh4_w6_22 :  std_logic;
signal bh4_w7_22 :  std_logic;
signal tile_23_X :  std_logic_vector(0 downto 0);
signal tile_23_Y :  std_logic_vector(7 downto 0);
signal tile_23_output :  std_logic_vector(7 downto 0);
signal tile_23_filtered_output :  unsigned(7-0 downto 0);
signal bh4_w0_23 :  std_logic;
signal bh4_w1_23 :  std_logic;
signal bh4_w2_23 :  std_logic;
signal bh4_w3_23 :  std_logic;
signal bh4_w4_23 :  std_logic;
signal bh4_w5_23 :  std_logic;
signal bh4_w6_23 :  std_logic;
signal bh4_w7_23 :  std_logic;
signal tile_24_X :  std_logic_vector(6 downto 0);
signal tile_24_Y :  std_logic_vector(0 downto 0);
signal tile_24_output :  std_logic_vector(6 downto 0);
signal tile_24_filtered_output :  unsigned(6-0 downto 0);
signal bh4_w0_24 :  std_logic;
signal bh4_w1_24 :  std_logic;
signal bh4_w2_24 :  std_logic;
signal bh4_w3_24 :  std_logic;
signal bh4_w4_24 :  std_logic;
signal bh4_w5_24 :  std_logic;
signal bh4_w6_24 :  std_logic;
signal tile_25_X :  std_logic_vector(0 downto 0);
signal tile_25_Y :  std_logic_vector(6 downto 0);
signal tile_25_output :  std_logic_vector(6 downto 0);
signal tile_25_filtered_output :  unsigned(6-0 downto 0);
signal bh4_w0_25 :  std_logic;
signal bh4_w1_25 :  std_logic;
signal bh4_w2_25 :  std_logic;
signal bh4_w3_25 :  std_logic;
signal bh4_w4_25 :  std_logic;
signal bh4_w5_25 :  std_logic;
signal bh4_w6_25 :  std_logic;
signal tile_26_X :  std_logic_vector(0 downto 0);
signal tile_26_Y :  std_logic_vector(5 downto 0);
signal tile_26_output :  std_logic_vector(5 downto 0);
signal tile_26_filtered_output :  unsigned(5-0 downto 0);
signal bh4_w0_26 :  std_logic;
signal bh4_w1_26 :  std_logic;
signal bh4_w2_26 :  std_logic;
signal bh4_w3_26 :  std_logic;
signal bh4_w4_26 :  std_logic;
signal bh4_w5_26 :  std_logic;
signal tile_27_X :  std_logic_vector(0 downto 0);
signal tile_27_Y :  std_logic_vector(4 downto 0);
signal tile_27_output :  std_logic_vector(4 downto 0);
signal tile_27_filtered_output :  unsigned(4-0 downto 0);
signal bh4_w0_27 :  std_logic;
signal bh4_w1_27 :  std_logic;
signal bh4_w2_27 :  std_logic;
signal bh4_w3_27 :  std_logic;
signal bh4_w4_27 :  std_logic;
signal tile_28_X :  std_logic_vector(4 downto 0);
signal tile_28_Y :  std_logic_vector(0 downto 0);
signal tile_28_output :  std_logic_vector(4 downto 0);
signal tile_28_filtered_output :  unsigned(4-0 downto 0);
signal bh4_w1_28 :  std_logic;
signal bh4_w2_28 :  std_logic;
signal bh4_w3_28 :  std_logic;
signal bh4_w4_28 :  std_logic;
signal bh4_w5_27 :  std_logic;
signal tile_29_X :  std_logic_vector(3 downto 0);
signal tile_29_Y :  std_logic_vector(0 downto 0);
signal tile_29_output :  std_logic_vector(3 downto 0);
signal tile_29_filtered_output :  unsigned(3-0 downto 0);
signal bh4_w1_29 :  std_logic;
signal bh4_w2_29 :  std_logic;
signal bh4_w3_29 :  std_logic;
signal bh4_w4_29 :  std_logic;
signal tile_30_X :  std_logic_vector(2 downto 0);
signal tile_30_Y :  std_logic_vector(18 downto 0);
signal tile_30_output :  std_logic_vector(21 downto 0);
signal tile_30_filtered_output :  unsigned(21-0 downto 0);
signal bh4_w17_4 :  std_logic;
signal bh4_w18_2 :  std_logic;
signal bh4_w19_1 :  std_logic;
signal bh4_w20_1 :  std_logic;
signal bh4_w21_1 :  std_logic;
signal bh4_w22_1 :  std_logic;
signal bh4_w23_1 :  std_logic;
signal bh4_w24_1 :  std_logic;
signal bh4_w25_1 :  std_logic;
signal bh4_w26_1 :  std_logic;
signal bh4_w27_1 :  std_logic;
signal bh4_w28_1 :  std_logic;
signal bh4_w29_1 :  std_logic;
signal bh4_w30_1 :  std_logic;
signal bh4_w31_1 :  std_logic;
signal bh4_w32_1 :  std_logic;
signal bh4_w33_1 :  std_logic;
signal bh4_w34_1 :  std_logic;
signal bh4_w35_1 :  std_logic;
signal bh4_w36_0 :  std_logic;
signal bh4_w37_0 :  std_logic;
signal bh4_w38_0 :  std_logic;
signal bh4_w0_28 :  std_logic;
signal bh4_w1_30 :  std_logic;
signal bh4_w2_30 :  std_logic;
signal bh4_w3_30 :  std_logic;
signal bh4_w4_30 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid70_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid70_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w0_29 :  std_logic;
signal bh4_w1_31 :  std_logic;
signal bh4_w2_31 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid70_Out0_copy71 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid72_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid72_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w0_30 :  std_logic;
signal bh4_w1_32 :  std_logic;
signal bh4_w2_32 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid72_Out0_copy73 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid74_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid74_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w0_31 :  std_logic;
signal bh4_w1_33 :  std_logic;
signal bh4_w2_33 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid74_Out0_copy75 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid76_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid76_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w0_32 :  std_logic;
signal bh4_w1_34 :  std_logic;
signal bh4_w2_34 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid76_Out0_copy77 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid80_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid80_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid80_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w0_33 :  std_logic;
signal bh4_w1_35 :  std_logic;
signal bh4_w2_35 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid80_Out0_copy81 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid82_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid82_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w1_36 :  std_logic;
signal bh4_w2_36 :  std_logic;
signal bh4_w3_31 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid82_Out0_copy83 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid84_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid84_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w1_37 :  std_logic;
signal bh4_w2_37 :  std_logic;
signal bh4_w3_32 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid84_Out0_copy85 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid86_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid86_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w1_38 :  std_logic;
signal bh4_w2_38 :  std_logic;
signal bh4_w3_33 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid86_Out0_copy87 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid88_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid88_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w1_39 :  std_logic;
signal bh4_w2_39 :  std_logic;
signal bh4_w3_34 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid88_Out0_copy89 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid90_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid90_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w1_40 :  std_logic;
signal bh4_w2_40 :  std_logic;
signal bh4_w3_35 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid90_Out0_copy91 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid92_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid92_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w2_41 :  std_logic;
signal bh4_w3_36 :  std_logic;
signal bh4_w4_31 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid92_Out0_copy93 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid94_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid94_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w2_42 :  std_logic;
signal bh4_w3_37 :  std_logic;
signal bh4_w4_32 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid94_Out0_copy95 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid96_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid96_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w2_43 :  std_logic;
signal bh4_w3_38 :  std_logic;
signal bh4_w4_33 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid96_Out0_copy97 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid98_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid98_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w2_44 :  std_logic;
signal bh4_w3_39 :  std_logic;
signal bh4_w4_34 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid98_Out0_copy99 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid100_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid100_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w2_45 :  std_logic;
signal bh4_w3_40 :  std_logic;
signal bh4_w4_35 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid100_Out0_copy101 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid102_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid102_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_41 :  std_logic;
signal bh4_w4_36 :  std_logic;
signal bh4_w5_28 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid102_Out0_copy103 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid104_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid104_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_42 :  std_logic;
signal bh4_w4_37 :  std_logic;
signal bh4_w5_29 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid104_Out0_copy105 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid106_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid106_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_43 :  std_logic;
signal bh4_w4_38 :  std_logic;
signal bh4_w5_30 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid106_Out0_copy107 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid108_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid108_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_44 :  std_logic;
signal bh4_w4_39 :  std_logic;
signal bh4_w5_31 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid108_Out0_copy109 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid110_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid110_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_45 :  std_logic;
signal bh4_w4_40 :  std_logic;
signal bh4_w5_32 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid110_Out0_copy111 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid112_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid112_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w4_41 :  std_logic;
signal bh4_w5_33 :  std_logic;
signal bh4_w6_26 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid112_Out0_copy113 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid114_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid114_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w4_42 :  std_logic;
signal bh4_w5_34 :  std_logic;
signal bh4_w6_27 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid114_Out0_copy115 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid116_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid116_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w4_43 :  std_logic;
signal bh4_w5_35 :  std_logic;
signal bh4_w6_28 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid116_Out0_copy117 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid118_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid118_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w4_44 :  std_logic;
signal bh4_w5_36 :  std_logic;
signal bh4_w6_29 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid118_Out0_copy119 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid120_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid120_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w4_45 :  std_logic;
signal bh4_w5_37 :  std_logic;
signal bh4_w6_30 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid120_Out0_copy121 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid122_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid122_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w5_38 :  std_logic;
signal bh4_w6_31 :  std_logic;
signal bh4_w7_24 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid122_Out0_copy123 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid124_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid124_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w5_39 :  std_logic;
signal bh4_w6_32 :  std_logic;
signal bh4_w7_25 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid124_Out0_copy125 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid126_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid126_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w5_40 :  std_logic;
signal bh4_w6_33 :  std_logic;
signal bh4_w7_26 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid126_Out0_copy127 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid128_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid128_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w5_41 :  std_logic;
signal bh4_w6_34 :  std_logic;
signal bh4_w7_27 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid128_Out0_copy129 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid130_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid130_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid130_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w5_42 :  std_logic;
signal bh4_w6_35 :  std_logic;
signal bh4_w7_28 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid130_Out0_copy131 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid132_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid132_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w6_36 :  std_logic;
signal bh4_w7_29 :  std_logic;
signal bh4_w8_22 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid132_Out0_copy133 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid134_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid134_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w6_37 :  std_logic;
signal bh4_w7_30 :  std_logic;
signal bh4_w8_23 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid134_Out0_copy135 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid136_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid136_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w6_38 :  std_logic;
signal bh4_w7_31 :  std_logic;
signal bh4_w8_24 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid136_Out0_copy137 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid138_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid138_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w6_39 :  std_logic;
signal bh4_w7_32 :  std_logic;
signal bh4_w8_25 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid138_Out0_copy139 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid140_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid140_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w7_33 :  std_logic;
signal bh4_w8_26 :  std_logic;
signal bh4_w9_20 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid140_Out0_copy141 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid142_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid142_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w7_34 :  std_logic;
signal bh4_w8_27 :  std_logic;
signal bh4_w9_21 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid142_Out0_copy143 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid144_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid144_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w7_35 :  std_logic;
signal bh4_w8_28 :  std_logic;
signal bh4_w9_22 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid144_Out0_copy145 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid146_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid146_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w7_36 :  std_logic;
signal bh4_w8_29 :  std_logic;
signal bh4_w9_23 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid146_Out0_copy147 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid148_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid148_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w8_30 :  std_logic;
signal bh4_w9_24 :  std_logic;
signal bh4_w10_18 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid148_Out0_copy149 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid150_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid150_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w8_31 :  std_logic;
signal bh4_w9_25 :  std_logic;
signal bh4_w10_19 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid150_Out0_copy151 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid152_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid152_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w8_32 :  std_logic;
signal bh4_w9_26 :  std_logic;
signal bh4_w10_20 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid152_Out0_copy153 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid154_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid154_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid154_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w8_33 :  std_logic;
signal bh4_w9_27 :  std_logic;
signal bh4_w10_21 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid154_Out0_copy155 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid156_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid156_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w9_28 :  std_logic;
signal bh4_w10_22 :  std_logic;
signal bh4_w11_16 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid156_Out0_copy157 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid158_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid158_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w9_29 :  std_logic;
signal bh4_w10_23 :  std_logic;
signal bh4_w11_17 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid158_Out0_copy159 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid160_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid160_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w9_30 :  std_logic;
signal bh4_w10_24 :  std_logic;
signal bh4_w11_18 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid160_Out0_copy161 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid162_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid162_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w10_25 :  std_logic;
signal bh4_w11_19 :  std_logic;
signal bh4_w12_14 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid162_Out0_copy163 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid164_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid164_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w10_26 :  std_logic;
signal bh4_w11_20 :  std_logic;
signal bh4_w12_15 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid164_Out0_copy165 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid166_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid166_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w10_27 :  std_logic;
signal bh4_w11_21 :  std_logic;
signal bh4_w12_16 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid166_Out0_copy167 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid168_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid168_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w11_22 :  std_logic;
signal bh4_w12_17 :  std_logic;
signal bh4_w13_12 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid168_Out0_copy169 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid170_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid170_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w11_23 :  std_logic;
signal bh4_w12_18 :  std_logic;
signal bh4_w13_13 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid170_Out0_copy171 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid172_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid172_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid172_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w11_24 :  std_logic;
signal bh4_w12_19 :  std_logic;
signal bh4_w13_14 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid172_Out0_copy173 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid174_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid174_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w12_20 :  std_logic;
signal bh4_w13_15 :  std_logic;
signal bh4_w14_10 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid174_Out0_copy175 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid176_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid176_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w12_21 :  std_logic;
signal bh4_w13_16 :  std_logic;
signal bh4_w14_11 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid176_Out0_copy177 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid178_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid178_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w13_17 :  std_logic;
signal bh4_w14_12 :  std_logic;
signal bh4_w15_8 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid178_Out0_copy179 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid180_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid180_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w13_18 :  std_logic;
signal bh4_w14_13 :  std_logic;
signal bh4_w15_9 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid180_Out0_copy181 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid182_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid182_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w14_14 :  std_logic;
signal bh4_w15_10 :  std_logic;
signal bh4_w16_6 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid182_Out0_copy183 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid184_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid184_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid184_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w14_15 :  std_logic;
signal bh4_w15_11 :  std_logic;
signal bh4_w16_7 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid184_Out0_copy185 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid186_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid186_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w15_12 :  std_logic;
signal bh4_w16_8 :  std_logic;
signal bh4_w17_5 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid186_Out0_copy187 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid188_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid188_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w16_9 :  std_logic;
signal bh4_w17_6 :  std_logic;
signal bh4_w18_3 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid188_Out0_copy189 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid190_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid190_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid190_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w17_7 :  std_logic;
signal bh4_w18_4 :  std_logic;
signal bh4_w19_2 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid190_Out0_copy191 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid194_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid194_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid194_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w18_5 :  std_logic;
signal bh4_w19_3 :  std_logic;
signal bh4_w20_2 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid194_Out0_copy195 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid196_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid196_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid196_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w20_3 :  std_logic;
signal bh4_w21_2 :  std_logic;
signal bh4_w22_2 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid196_Out0_copy197 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid198_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid198_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid198_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w22_3 :  std_logic;
signal bh4_w23_2 :  std_logic;
signal bh4_w24_2 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid198_Out0_copy199 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid200_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid200_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid200_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w24_3 :  std_logic;
signal bh4_w25_2 :  std_logic;
signal bh4_w26_2 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid200_Out0_copy201 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid202_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid202_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid202_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w26_3 :  std_logic;
signal bh4_w27_2 :  std_logic;
signal bh4_w28_2 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid202_Out0_copy203 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid204_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid204_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid204_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w28_3 :  std_logic;
signal bh4_w29_2 :  std_logic;
signal bh4_w30_2 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid204_Out0_copy205 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid206_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid206_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid206_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w30_3 :  std_logic;
signal bh4_w31_2 :  std_logic;
signal bh4_w32_2 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid206_Out0_copy207 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid208_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid208_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid208_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w32_3 :  std_logic;
signal bh4_w33_2 :  std_logic;
signal bh4_w34_2 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid208_Out0_copy209 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid210_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid210_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid210_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w34_3 :  std_logic;
signal bh4_w35_2 :  std_logic;
signal bh4_w36_1 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid210_Out0_copy211 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid212_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid212_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w0_34 :  std_logic;
signal bh4_w1_41 :  std_logic;
signal bh4_w2_46 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid212_Out0_copy213 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid214_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid214_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w1_42 :  std_logic;
signal bh4_w2_47 :  std_logic;
signal bh4_w3_46 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid214_Out0_copy215 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid216_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid216_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid216_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w1_43 :  std_logic;
signal bh4_w2_48 :  std_logic;
signal bh4_w3_47 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid216_Out0_copy217 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid218_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid218_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w2_49 :  std_logic;
signal bh4_w3_48 :  std_logic;
signal bh4_w4_46 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid218_Out0_copy219 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid220_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid220_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w2_50 :  std_logic;
signal bh4_w3_49 :  std_logic;
signal bh4_w4_47 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid220_Out0_copy221 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid224_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid224_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w2_51 :  std_logic;
signal bh4_w3_50 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid224_Out0_copy225 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid226_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid226_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_51 :  std_logic;
signal bh4_w4_48 :  std_logic;
signal bh4_w5_43 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid226_Out0_copy227 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid228_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid228_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_52 :  std_logic;
signal bh4_w4_49 :  std_logic;
signal bh4_w5_44 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid228_Out0_copy229 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid230_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid230_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid230_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_53 :  std_logic;
signal bh4_w4_50 :  std_logic;
signal bh4_w5_45 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid230_Out0_copy231 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid232_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid232_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w4_51 :  std_logic;
signal bh4_w5_46 :  std_logic;
signal bh4_w6_40 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid232_Out0_copy233 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid234_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid234_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w4_52 :  std_logic;
signal bh4_w5_47 :  std_logic;
signal bh4_w6_41 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid234_Out0_copy235 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid236_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid236_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid236_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w4_53 :  std_logic;
signal bh4_w5_48 :  std_logic;
signal bh4_w6_42 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid236_Out0_copy237 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid238_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid238_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w5_49 :  std_logic;
signal bh4_w6_43 :  std_logic;
signal bh4_w7_37 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid238_Out0_copy239 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid240_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid240_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w5_50 :  std_logic;
signal bh4_w6_44 :  std_logic;
signal bh4_w7_38 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid240_Out0_copy241 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid242_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid242_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w6_45 :  std_logic;
signal bh4_w7_39 :  std_logic;
signal bh4_w8_34 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid242_Out0_copy243 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid244_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid244_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w6_46 :  std_logic;
signal bh4_w7_40 :  std_logic;
signal bh4_w8_35 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid244_Out0_copy245 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid246_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid246_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w6_47 :  std_logic;
signal bh4_w7_41 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid246_Out0_copy247 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid248_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid248_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w7_42 :  std_logic;
signal bh4_w8_36 :  std_logic;
signal bh4_w9_31 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid248_Out0_copy249 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid250_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid250_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w7_43 :  std_logic;
signal bh4_w8_37 :  std_logic;
signal bh4_w9_32 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid250_Out0_copy251 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid252_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid252_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w8_38 :  std_logic;
signal bh4_w9_33 :  std_logic;
signal bh4_w10_28 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid252_Out0_copy253 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid254_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid254_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w8_39 :  std_logic;
signal bh4_w9_34 :  std_logic;
signal bh4_w10_29 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid254_Out0_copy255 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid256_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid256_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w9_35 :  std_logic;
signal bh4_w10_30 :  std_logic;
signal bh4_w11_25 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid256_Out0_copy257 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid258_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid258_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w9_36 :  std_logic;
signal bh4_w10_31 :  std_logic;
signal bh4_w11_26 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid258_Out0_copy259 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid260_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid260_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w10_32 :  std_logic;
signal bh4_w11_27 :  std_logic;
signal bh4_w12_22 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid260_Out0_copy261 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid262_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid262_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid262_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w10_33 :  std_logic;
signal bh4_w11_28 :  std_logic;
signal bh4_w12_23 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid262_Out0_copy263 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid264_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid264_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w11_29 :  std_logic;
signal bh4_w12_24 :  std_logic;
signal bh4_w13_19 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid264_Out0_copy265 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid266_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid266_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w11_30 :  std_logic;
signal bh4_w12_25 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid266_Out0_copy267 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid268_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid268_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w12_26 :  std_logic;
signal bh4_w13_20 :  std_logic;
signal bh4_w14_16 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid268_Out0_copy269 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid270_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid270_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w12_27 :  std_logic;
signal bh4_w13_21 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid270_Out0_copy271 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid272_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid272_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w13_22 :  std_logic;
signal bh4_w14_17 :  std_logic;
signal bh4_w15_13 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid272_Out0_copy273 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid274_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid274_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w14_18 :  std_logic;
signal bh4_w15_14 :  std_logic;
signal bh4_w16_10 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid274_Out0_copy275 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid276_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid276_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w15_15 :  std_logic;
signal bh4_w16_11 :  std_logic;
signal bh4_w17_8 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid276_Out0_copy277 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid278_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid278_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid278_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w16_12 :  std_logic;
signal bh4_w17_9 :  std_logic;
signal bh4_w18_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid278_Out0_copy279 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid280_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid280_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid280_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w17_10 :  std_logic;
signal bh4_w18_7 :  std_logic;
signal bh4_w19_4 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid280_Out0_copy281 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid282_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid282_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid282_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w19_5 :  std_logic;
signal bh4_w20_4 :  std_logic;
signal bh4_w21_3 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid282_Out0_copy283 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid284_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid284_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid284_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w22_4 :  std_logic;
signal bh4_w23_3 :  std_logic;
signal bh4_w24_4 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid284_Out0_copy285 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid286_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid286_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid286_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w24_5 :  std_logic;
signal bh4_w25_3 :  std_logic;
signal bh4_w26_4 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid286_Out0_copy287 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid288_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid288_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid288_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w26_5 :  std_logic;
signal bh4_w27_3 :  std_logic;
signal bh4_w28_4 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid288_Out0_copy289 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid290_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid290_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid290_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w28_5 :  std_logic;
signal bh4_w29_3 :  std_logic;
signal bh4_w30_4 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid290_Out0_copy291 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid292_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid292_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid292_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w30_5 :  std_logic;
signal bh4_w31_3 :  std_logic;
signal bh4_w32_4 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid292_Out0_copy293 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid294_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid294_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid294_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w32_5 :  std_logic;
signal bh4_w33_3 :  std_logic;
signal bh4_w34_4 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid294_Out0_copy295 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid296_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid296_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid296_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w34_5 :  std_logic;
signal bh4_w35_3 :  std_logic;
signal bh4_w36_2 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid296_Out0_copy297 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid298_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid298_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid298_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w36_3 :  std_logic;
signal bh4_w37_1 :  std_logic;
signal bh4_w38_1 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid298_Out0_copy299 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid300_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid300_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w1_44 :  std_logic;
signal bh4_w2_52 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid300_Out0_copy301 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid302_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid302_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w2_53 :  std_logic;
signal bh4_w3_54 :  std_logic;
signal bh4_w4_54 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid302_Out0_copy303 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid304_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid304_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_55 :  std_logic;
signal bh4_w4_55 :  std_logic;
signal bh4_w5_51 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid304_Out0_copy305 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid306_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid306_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid306_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_56 :  std_logic;
signal bh4_w4_56 :  std_logic;
signal bh4_w5_52 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid306_Out0_copy307 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid308_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid308_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w4_57 :  std_logic;
signal bh4_w5_53 :  std_logic;
signal bh4_w6_48 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid308_Out0_copy309 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid310_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid310_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w5_54 :  std_logic;
signal bh4_w6_49 :  std_logic;
signal bh4_w7_44 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid310_Out0_copy311 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid312_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid312_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid312_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w5_55 :  std_logic;
signal bh4_w6_50 :  std_logic;
signal bh4_w7_45 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid312_Out0_copy313 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid314_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid314_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w6_51 :  std_logic;
signal bh4_w7_46 :  std_logic;
signal bh4_w8_40 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid314_Out0_copy315 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid316_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid316_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w7_47 :  std_logic;
signal bh4_w8_41 :  std_logic;
signal bh4_w9_37 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid316_Out0_copy317 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid318_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid318_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w7_48 :  std_logic;
signal bh4_w8_42 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid318_Out0_copy319 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid320_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid320_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w8_43 :  std_logic;
signal bh4_w9_38 :  std_logic;
signal bh4_w10_34 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid320_Out0_copy321 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid322_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid322_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w9_39 :  std_logic;
signal bh4_w10_35 :  std_logic;
signal bh4_w11_31 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid322_Out0_copy323 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid324_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid324_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w10_36 :  std_logic;
signal bh4_w11_32 :  std_logic;
signal bh4_w12_28 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid324_Out0_copy325 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid326_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid326_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w11_33 :  std_logic;
signal bh4_w12_29 :  std_logic;
signal bh4_w13_23 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid326_Out0_copy327 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid328_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F125_uid69_bh4_uid328_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w12_30 :  std_logic;
signal bh4_w13_24 :  std_logic;
signal bh4_w14_19 :  std_logic;
signal Compressor_6_3_F125_uid69_bh4_uid328_Out0_copy329 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid330_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid330_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid330_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w13_25 :  std_logic;
signal bh4_w14_20 :  std_logic;
signal bh4_w15_16 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid330_Out0_copy331 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid332_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid332_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid332_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w13_26 :  std_logic;
signal bh4_w14_21 :  std_logic;
signal bh4_w15_17 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid332_Out0_copy333 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid334_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid334_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid334_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w15_18 :  std_logic;
signal bh4_w16_13 :  std_logic;
signal bh4_w17_11 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid334_Out0_copy335 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid336_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid336_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid336_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w17_12 :  std_logic;
signal bh4_w18_8 :  std_logic;
signal bh4_w19_6 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid336_Out0_copy337 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid338_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid338_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid338_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w19_7 :  std_logic;
signal bh4_w20_5 :  std_logic;
signal bh4_w21_4 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid338_Out0_copy339 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid340_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid340_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid340_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w21_5 :  std_logic;
signal bh4_w22_5 :  std_logic;
signal bh4_w23_4 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid340_Out0_copy341 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid342_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid342_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid342_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w24_6 :  std_logic;
signal bh4_w25_4 :  std_logic;
signal bh4_w26_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid342_Out0_copy343 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid344_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid344_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid344_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w26_7 :  std_logic;
signal bh4_w27_4 :  std_logic;
signal bh4_w28_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid344_Out0_copy345 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid346_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid346_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid346_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w28_7 :  std_logic;
signal bh4_w29_4 :  std_logic;
signal bh4_w30_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid346_Out0_copy347 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid348_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid348_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid348_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w30_7 :  std_logic;
signal bh4_w31_4 :  std_logic;
signal bh4_w32_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid348_Out0_copy349 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid350_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid350_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid350_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w32_7 :  std_logic;
signal bh4_w33_4 :  std_logic;
signal bh4_w34_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid350_Out0_copy351 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid352_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid352_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid352_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w34_7 :  std_logic;
signal bh4_w35_4 :  std_logic;
signal bh4_w36_4 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid352_Out0_copy353 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid354_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid354_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid354_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w36_5 :  std_logic;
signal bh4_w37_2 :  std_logic;
signal bh4_w38_2 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid354_Out0_copy355 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid356_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid356_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w38_3 :  std_logic;
signal bh4_w39_0 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid356_Out0_copy357 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid358_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid358_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid358_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w1_45 :  std_logic;
signal bh4_w2_54 :  std_logic;
signal bh4_w3_57 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid358_Out0_copy359 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid360_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid360_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w3_58 :  std_logic;
signal bh4_w4_58 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid360_Out0_copy361 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid362_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid362_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid362_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w4_59 :  std_logic;
signal bh4_w5_56 :  std_logic;
signal bh4_w6_52 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid362_Out0_copy363 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid364_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid364_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid364_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w5_57 :  std_logic;
signal bh4_w6_53 :  std_logic;
signal bh4_w7_49 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid364_Out0_copy365 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid366_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid366_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w6_54 :  std_logic;
signal bh4_w7_50 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid366_Out0_copy367 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid368_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid368_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid368_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w7_51 :  std_logic;
signal bh4_w8_44 :  std_logic;
signal bh4_w9_40 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid368_Out0_copy369 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid370_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid370_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid370_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w8_45 :  std_logic;
signal bh4_w9_41 :  std_logic;
signal bh4_w10_37 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid370_Out0_copy371 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid372_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid372_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid372_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w10_38 :  std_logic;
signal bh4_w11_34 :  std_logic;
signal bh4_w12_31 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid372_Out0_copy373 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid374_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid374_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w12_32 :  std_logic;
signal bh4_w13_27 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid374_Out0_copy375 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid376_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid376_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid376_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w13_28 :  std_logic;
signal bh4_w14_22 :  std_logic;
signal bh4_w15_19 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid376_Out0_copy377 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid378_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid378_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w14_23 :  std_logic;
signal bh4_w15_20 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid378_Out0_copy379 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid380_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid380_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid380_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w15_21 :  std_logic;
signal bh4_w16_14 :  std_logic;
signal bh4_w17_13 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid380_Out0_copy381 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid382_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid382_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid382_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w17_14 :  std_logic;
signal bh4_w18_9 :  std_logic;
signal bh4_w19_8 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid382_Out0_copy383 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid384_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid384_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid384_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w19_9 :  std_logic;
signal bh4_w20_6 :  std_logic;
signal bh4_w21_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid384_Out0_copy385 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid386_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid386_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid386_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w21_7 :  std_logic;
signal bh4_w22_6 :  std_logic;
signal bh4_w23_5 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid386_Out0_copy387 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid388_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid388_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid388_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w23_6 :  std_logic;
signal bh4_w24_7 :  std_logic;
signal bh4_w25_5 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid388_Out0_copy389 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid390_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid390_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid390_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w26_8 :  std_logic;
signal bh4_w27_5 :  std_logic;
signal bh4_w28_8 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid390_Out0_copy391 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid392_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid392_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid392_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w28_9 :  std_logic;
signal bh4_w29_5 :  std_logic;
signal bh4_w30_8 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid392_Out0_copy393 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid394_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid394_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid394_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w30_9 :  std_logic;
signal bh4_w31_5 :  std_logic;
signal bh4_w32_8 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid394_Out0_copy395 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid396_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid396_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid396_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w32_9 :  std_logic;
signal bh4_w33_5 :  std_logic;
signal bh4_w34_8 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid396_Out0_copy397 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid398_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid398_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid398_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w34_9 :  std_logic;
signal bh4_w35_5 :  std_logic;
signal bh4_w36_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid398_Out0_copy399 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid400_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid400_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid400_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w36_7 :  std_logic;
signal bh4_w37_3 :  std_logic;
signal bh4_w38_4 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid400_Out0_copy401 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid402_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid402_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid402_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w38_5 :  std_logic;
signal bh4_w39_1 :  std_logic;
signal bh4_w40_0 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid402_Out0_copy403 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid404_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid404_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid404_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w3_59 :  std_logic;
signal bh4_w4_60 :  std_logic;
signal bh4_w5_58 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid404_Out0_copy405 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid406_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid406_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w5_59 :  std_logic;
signal bh4_w6_55 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid406_Out0_copy407 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid408_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid408_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w6_56 :  std_logic;
signal bh4_w7_52 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid408_Out0_copy409 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid410_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid410_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid410_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w7_53 :  std_logic;
signal bh4_w8_46 :  std_logic;
signal bh4_w9_42 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid410_Out0_copy411 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid412_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid412_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid412_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w9_43 :  std_logic;
signal bh4_w10_39 :  std_logic;
signal bh4_w11_35 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid412_Out0_copy413 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid414_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid414_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid414_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w11_36 :  std_logic;
signal bh4_w12_33 :  std_logic;
signal bh4_w13_29 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid414_Out0_copy415 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid416_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid416_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F125_uid193_bh4_uid416_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w13_30 :  std_logic;
signal bh4_w14_24 :  std_logic;
signal bh4_w15_22 :  std_logic;
signal Compressor_23_3_F125_uid193_bh4_uid416_Out0_copy417 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid418_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F125_uid223_bh4_uid418_Out0 :  std_logic_vector(1 downto 0);
signal bh4_w15_23 :  std_logic;
signal bh4_w16_15 :  std_logic;
signal Compressor_3_2_F125_uid223_bh4_uid418_Out0_copy419 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid420_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid420_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid420_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w17_15 :  std_logic;
signal bh4_w18_10 :  std_logic;
signal bh4_w19_10 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid420_Out0_copy421 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid422_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid422_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid422_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w19_11 :  std_logic;
signal bh4_w20_7 :  std_logic;
signal bh4_w21_8 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid422_Out0_copy423 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid424_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid424_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid424_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w21_9 :  std_logic;
signal bh4_w22_7 :  std_logic;
signal bh4_w23_7 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid424_Out0_copy425 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid426_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid426_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid426_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w23_8 :  std_logic;
signal bh4_w24_8 :  std_logic;
signal bh4_w25_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid426_Out0_copy427 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid428_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid428_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid428_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w25_7 :  std_logic;
signal bh4_w26_9 :  std_logic;
signal bh4_w27_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid428_Out0_copy429 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid430_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid430_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid430_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w28_10 :  std_logic;
signal bh4_w29_6 :  std_logic;
signal bh4_w30_10 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid430_Out0_copy431 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid432_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid432_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid432_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w30_11 :  std_logic;
signal bh4_w31_6 :  std_logic;
signal bh4_w32_10 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid432_Out0_copy433 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid434_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid434_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid434_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w32_11 :  std_logic;
signal bh4_w33_6 :  std_logic;
signal bh4_w34_10 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid434_Out0_copy435 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid436_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid436_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid436_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w34_11 :  std_logic;
signal bh4_w35_6 :  std_logic;
signal bh4_w36_8 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid436_Out0_copy437 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid438_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid438_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid438_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w36_9 :  std_logic;
signal bh4_w37_4 :  std_logic;
signal bh4_w38_6 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid438_Out0_copy439 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid440_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid440_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F125_uid79_bh4_uid440_Out0 :  std_logic_vector(2 downto 0);
signal bh4_w38_7 :  std_logic;
signal bh4_w39_2 :  std_logic;
signal bh4_w40_1 :  std_logic;
signal Compressor_14_3_F125_uid79_bh4_uid440_Out0_copy441 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh4_4 :  std_logic_vector(4 downto 0);
signal bitheapFinalAdd_bh4_In0 :  std_logic_vector(63 downto 0);
signal bitheapFinalAdd_bh4_In1 :  std_logic_vector(63 downto 0);
signal bitheapFinalAdd_bh4_Cin :  std_logic;
signal bitheapFinalAdd_bh4_Out :  std_logic_vector(63 downto 0);
signal bitheapResult_bh4 :  std_logic_vector(67 downto 0);
begin
   XX_m3 <= X ;
   YY_m3 <= Y ;
   tile_0_X <= X(30 downto 14);
   tile_0_Y <= Y(33 downto 15);
   tile_0_mult: DSPBlock_17x19_F125_uid6
      port map ( clk  => clk,
                 X => tile_0_X,
                 Y => tile_0_Y,
                 R => tile_0_output);

   tile_0_filtered_output <= unsigned(tile_0_output(35 downto 0));
   bh4_w0_0 <= tile_0_filtered_output(0);
   bh4_w1_0 <= tile_0_filtered_output(1);
   bh4_w2_0 <= tile_0_filtered_output(2);
   bh4_w3_0 <= tile_0_filtered_output(3);
   bh4_w4_0 <= tile_0_filtered_output(4);
   bh4_w5_0 <= tile_0_filtered_output(5);
   bh4_w6_0 <= tile_0_filtered_output(6);
   bh4_w7_0 <= tile_0_filtered_output(7);
   bh4_w8_0 <= tile_0_filtered_output(8);
   bh4_w9_0 <= tile_0_filtered_output(9);
   bh4_w10_0 <= tile_0_filtered_output(10);
   bh4_w11_0 <= tile_0_filtered_output(11);
   bh4_w12_0 <= tile_0_filtered_output(12);
   bh4_w13_0 <= tile_0_filtered_output(13);
   bh4_w14_0 <= tile_0_filtered_output(14);
   bh4_w15_0 <= tile_0_filtered_output(15);
   bh4_w16_0 <= tile_0_filtered_output(16);
   bh4_w17_0 <= tile_0_filtered_output(17);
   bh4_w18_0 <= tile_0_filtered_output(18);
   bh4_w19_0 <= tile_0_filtered_output(19);
   bh4_w20_0 <= tile_0_filtered_output(20);
   bh4_w21_0 <= tile_0_filtered_output(21);
   bh4_w22_0 <= tile_0_filtered_output(22);
   bh4_w23_0 <= tile_0_filtered_output(23);
   bh4_w24_0 <= tile_0_filtered_output(24);
   bh4_w25_0 <= tile_0_filtered_output(25);
   bh4_w26_0 <= tile_0_filtered_output(26);
   bh4_w27_0 <= tile_0_filtered_output(27);
   bh4_w28_0 <= tile_0_filtered_output(28);
   bh4_w29_0 <= tile_0_filtered_output(29);
   bh4_w30_0 <= tile_0_filtered_output(30);
   bh4_w31_0 <= tile_0_filtered_output(31);
   bh4_w32_0 <= tile_0_filtered_output(32);
   bh4_w33_0 <= tile_0_filtered_output(33);
   bh4_w34_0 <= tile_0_filtered_output(34);
   bh4_w35_0 <= tile_0_filtered_output(35);
   tile_1_X <= X(33 downto 15);
   tile_1_Y <= Y(14 downto 14);
   tile_1_mult: DSPBlock_19x1_F125_uid8
      port map ( clk  => clk,
                 X => tile_1_X,
                 Y => tile_1_Y,
                 R => tile_1_output);

   tile_1_filtered_output <= unsigned(tile_1_output(18 downto 0));
   bh4_w0_1 <= tile_1_filtered_output(0);
   bh4_w1_1 <= tile_1_filtered_output(1);
   bh4_w2_1 <= tile_1_filtered_output(2);
   bh4_w3_1 <= tile_1_filtered_output(3);
   bh4_w4_1 <= tile_1_filtered_output(4);
   bh4_w5_1 <= tile_1_filtered_output(5);
   bh4_w6_1 <= tile_1_filtered_output(6);
   bh4_w7_1 <= tile_1_filtered_output(7);
   bh4_w8_1 <= tile_1_filtered_output(8);
   bh4_w9_1 <= tile_1_filtered_output(9);
   bh4_w10_1 <= tile_1_filtered_output(10);
   bh4_w11_1 <= tile_1_filtered_output(11);
   bh4_w12_1 <= tile_1_filtered_output(12);
   bh4_w13_1 <= tile_1_filtered_output(13);
   bh4_w14_1 <= tile_1_filtered_output(14);
   bh4_w15_1 <= tile_1_filtered_output(15);
   bh4_w16_1 <= tile_1_filtered_output(16);
   bh4_w17_1 <= tile_1_filtered_output(17);
   bh4_w18_1 <= tile_1_filtered_output(18);
   tile_2_X <= X(33 downto 16);
   tile_2_Y <= Y(13 downto 13);
   tile_2_mult: DSPBlock_18x1_F125_uid10
      port map ( clk  => clk,
                 X => tile_2_X,
                 Y => tile_2_Y,
                 R => tile_2_output);

   tile_2_filtered_output <= unsigned(tile_2_output(17 downto 0));
   bh4_w0_2 <= tile_2_filtered_output(0);
   bh4_w1_2 <= tile_2_filtered_output(1);
   bh4_w2_2 <= tile_2_filtered_output(2);
   bh4_w3_2 <= tile_2_filtered_output(3);
   bh4_w4_2 <= tile_2_filtered_output(4);
   bh4_w5_2 <= tile_2_filtered_output(5);
   bh4_w6_2 <= tile_2_filtered_output(6);
   bh4_w7_2 <= tile_2_filtered_output(7);
   bh4_w8_2 <= tile_2_filtered_output(8);
   bh4_w9_2 <= tile_2_filtered_output(9);
   bh4_w10_2 <= tile_2_filtered_output(10);
   bh4_w11_2 <= tile_2_filtered_output(11);
   bh4_w12_2 <= tile_2_filtered_output(12);
   bh4_w13_2 <= tile_2_filtered_output(13);
   bh4_w14_2 <= tile_2_filtered_output(14);
   bh4_w15_2 <= tile_2_filtered_output(15);
   bh4_w16_2 <= tile_2_filtered_output(16);
   bh4_w17_2 <= tile_2_filtered_output(17);
   tile_3_X <= X(13 downto 13);
   tile_3_Y <= Y(33 downto 16);
   tile_3_mult: DSPBlock_1x18_F125_uid12
      port map ( clk  => clk,
                 X => tile_3_X,
                 Y => tile_3_Y,
                 R => tile_3_output);

   tile_3_filtered_output <= unsigned(tile_3_output(17 downto 0));
   bh4_w0_3 <= tile_3_filtered_output(0);
   bh4_w1_3 <= tile_3_filtered_output(1);
   bh4_w2_3 <= tile_3_filtered_output(2);
   bh4_w3_3 <= tile_3_filtered_output(3);
   bh4_w4_3 <= tile_3_filtered_output(4);
   bh4_w5_3 <= tile_3_filtered_output(5);
   bh4_w6_3 <= tile_3_filtered_output(6);
   bh4_w7_3 <= tile_3_filtered_output(7);
   bh4_w8_3 <= tile_3_filtered_output(8);
   bh4_w9_3 <= tile_3_filtered_output(9);
   bh4_w10_3 <= tile_3_filtered_output(10);
   bh4_w11_3 <= tile_3_filtered_output(11);
   bh4_w12_3 <= tile_3_filtered_output(12);
   bh4_w13_3 <= tile_3_filtered_output(13);
   bh4_w14_3 <= tile_3_filtered_output(14);
   bh4_w15_3 <= tile_3_filtered_output(15);
   bh4_w16_3 <= tile_3_filtered_output(16);
   bh4_w17_3 <= tile_3_filtered_output(17);
   tile_4_X <= X(12 downto 12);
   tile_4_Y <= Y(33 downto 17);
   tile_4_mult: DSPBlock_1x17_F125_uid14
      port map ( clk  => clk,
                 X => tile_4_X,
                 Y => tile_4_Y,
                 R => tile_4_output);

   tile_4_filtered_output <= unsigned(tile_4_output(16 downto 0));
   bh4_w0_4 <= tile_4_filtered_output(0);
   bh4_w1_4 <= tile_4_filtered_output(1);
   bh4_w2_4 <= tile_4_filtered_output(2);
   bh4_w3_4 <= tile_4_filtered_output(3);
   bh4_w4_4 <= tile_4_filtered_output(4);
   bh4_w5_4 <= tile_4_filtered_output(5);
   bh4_w6_4 <= tile_4_filtered_output(6);
   bh4_w7_4 <= tile_4_filtered_output(7);
   bh4_w8_4 <= tile_4_filtered_output(8);
   bh4_w9_4 <= tile_4_filtered_output(9);
   bh4_w10_4 <= tile_4_filtered_output(10);
   bh4_w11_4 <= tile_4_filtered_output(11);
   bh4_w12_4 <= tile_4_filtered_output(12);
   bh4_w13_4 <= tile_4_filtered_output(13);
   bh4_w14_4 <= tile_4_filtered_output(14);
   bh4_w15_4 <= tile_4_filtered_output(15);
   bh4_w16_4 <= tile_4_filtered_output(16);
   tile_5_X <= X(33 downto 17);
   tile_5_Y <= Y(12 downto 12);
   tile_5_mult: DSPBlock_17x1_F125_uid16
      port map ( clk  => clk,
                 X => tile_5_X,
                 Y => tile_5_Y,
                 R => tile_5_output);

   tile_5_filtered_output <= unsigned(tile_5_output(16 downto 0));
   bh4_w0_5 <= tile_5_filtered_output(0);
   bh4_w1_5 <= tile_5_filtered_output(1);
   bh4_w2_5 <= tile_5_filtered_output(2);
   bh4_w3_5 <= tile_5_filtered_output(3);
   bh4_w4_5 <= tile_5_filtered_output(4);
   bh4_w5_5 <= tile_5_filtered_output(5);
   bh4_w6_5 <= tile_5_filtered_output(6);
   bh4_w7_5 <= tile_5_filtered_output(7);
   bh4_w8_5 <= tile_5_filtered_output(8);
   bh4_w9_5 <= tile_5_filtered_output(9);
   bh4_w10_5 <= tile_5_filtered_output(10);
   bh4_w11_5 <= tile_5_filtered_output(11);
   bh4_w12_5 <= tile_5_filtered_output(12);
   bh4_w13_5 <= tile_5_filtered_output(13);
   bh4_w14_5 <= tile_5_filtered_output(14);
   bh4_w15_5 <= tile_5_filtered_output(15);
   bh4_w16_5 <= tile_5_filtered_output(16);
   tile_6_X <= X(33 downto 18);
   tile_6_Y <= Y(11 downto 11);
   tile_6_mult: DSPBlock_16x1_F125_uid18
      port map ( clk  => clk,
                 X => tile_6_X,
                 Y => tile_6_Y,
                 R => tile_6_output);

   tile_6_filtered_output <= unsigned(tile_6_output(15 downto 0));
   bh4_w0_6 <= tile_6_filtered_output(0);
   bh4_w1_6 <= tile_6_filtered_output(1);
   bh4_w2_6 <= tile_6_filtered_output(2);
   bh4_w3_6 <= tile_6_filtered_output(3);
   bh4_w4_6 <= tile_6_filtered_output(4);
   bh4_w5_6 <= tile_6_filtered_output(5);
   bh4_w6_6 <= tile_6_filtered_output(6);
   bh4_w7_6 <= tile_6_filtered_output(7);
   bh4_w8_6 <= tile_6_filtered_output(8);
   bh4_w9_6 <= tile_6_filtered_output(9);
   bh4_w10_6 <= tile_6_filtered_output(10);
   bh4_w11_6 <= tile_6_filtered_output(11);
   bh4_w12_6 <= tile_6_filtered_output(12);
   bh4_w13_6 <= tile_6_filtered_output(13);
   bh4_w14_6 <= tile_6_filtered_output(14);
   bh4_w15_6 <= tile_6_filtered_output(15);
   tile_7_X <= X(11 downto 11);
   tile_7_Y <= Y(33 downto 18);
   tile_7_mult: DSPBlock_1x16_F125_uid20
      port map ( clk  => clk,
                 X => tile_7_X,
                 Y => tile_7_Y,
                 R => tile_7_output);

   tile_7_filtered_output <= unsigned(tile_7_output(15 downto 0));
   bh4_w0_7 <= tile_7_filtered_output(0);
   bh4_w1_7 <= tile_7_filtered_output(1);
   bh4_w2_7 <= tile_7_filtered_output(2);
   bh4_w3_7 <= tile_7_filtered_output(3);
   bh4_w4_7 <= tile_7_filtered_output(4);
   bh4_w5_7 <= tile_7_filtered_output(5);
   bh4_w6_7 <= tile_7_filtered_output(6);
   bh4_w7_7 <= tile_7_filtered_output(7);
   bh4_w8_7 <= tile_7_filtered_output(8);
   bh4_w9_7 <= tile_7_filtered_output(9);
   bh4_w10_7 <= tile_7_filtered_output(10);
   bh4_w11_7 <= tile_7_filtered_output(11);
   bh4_w12_7 <= tile_7_filtered_output(12);
   bh4_w13_7 <= tile_7_filtered_output(13);
   bh4_w14_7 <= tile_7_filtered_output(14);
   bh4_w15_7 <= tile_7_filtered_output(15);
   tile_8_X <= X(10 downto 10);
   tile_8_Y <= Y(33 downto 19);
   tile_8_mult: DSPBlock_1x15_F125_uid22
      port map ( clk  => clk,
                 X => tile_8_X,
                 Y => tile_8_Y,
                 R => tile_8_output);

   tile_8_filtered_output <= unsigned(tile_8_output(14 downto 0));
   bh4_w0_8 <= tile_8_filtered_output(0);
   bh4_w1_8 <= tile_8_filtered_output(1);
   bh4_w2_8 <= tile_8_filtered_output(2);
   bh4_w3_8 <= tile_8_filtered_output(3);
   bh4_w4_8 <= tile_8_filtered_output(4);
   bh4_w5_8 <= tile_8_filtered_output(5);
   bh4_w6_8 <= tile_8_filtered_output(6);
   bh4_w7_8 <= tile_8_filtered_output(7);
   bh4_w8_8 <= tile_8_filtered_output(8);
   bh4_w9_8 <= tile_8_filtered_output(9);
   bh4_w10_8 <= tile_8_filtered_output(10);
   bh4_w11_8 <= tile_8_filtered_output(11);
   bh4_w12_8 <= tile_8_filtered_output(12);
   bh4_w13_8 <= tile_8_filtered_output(13);
   bh4_w14_8 <= tile_8_filtered_output(14);
   tile_9_X <= X(33 downto 19);
   tile_9_Y <= Y(10 downto 10);
   tile_9_mult: DSPBlock_15x1_F125_uid24
      port map ( clk  => clk,
                 X => tile_9_X,
                 Y => tile_9_Y,
                 R => tile_9_output);

   tile_9_filtered_output <= unsigned(tile_9_output(14 downto 0));
   bh4_w0_9 <= tile_9_filtered_output(0);
   bh4_w1_9 <= tile_9_filtered_output(1);
   bh4_w2_9 <= tile_9_filtered_output(2);
   bh4_w3_9 <= tile_9_filtered_output(3);
   bh4_w4_9 <= tile_9_filtered_output(4);
   bh4_w5_9 <= tile_9_filtered_output(5);
   bh4_w6_9 <= tile_9_filtered_output(6);
   bh4_w7_9 <= tile_9_filtered_output(7);
   bh4_w8_9 <= tile_9_filtered_output(8);
   bh4_w9_9 <= tile_9_filtered_output(9);
   bh4_w10_9 <= tile_9_filtered_output(10);
   bh4_w11_9 <= tile_9_filtered_output(11);
   bh4_w12_9 <= tile_9_filtered_output(12);
   bh4_w13_9 <= tile_9_filtered_output(13);
   bh4_w14_9 <= tile_9_filtered_output(14);
   tile_10_X <= X(33 downto 20);
   tile_10_Y <= Y(9 downto 9);
   tile_10_mult: DSPBlock_14x1_F125_uid26
      port map ( clk  => clk,
                 X => tile_10_X,
                 Y => tile_10_Y,
                 R => tile_10_output);

   tile_10_filtered_output <= unsigned(tile_10_output(13 downto 0));
   bh4_w0_10 <= tile_10_filtered_output(0);
   bh4_w1_10 <= tile_10_filtered_output(1);
   bh4_w2_10 <= tile_10_filtered_output(2);
   bh4_w3_10 <= tile_10_filtered_output(3);
   bh4_w4_10 <= tile_10_filtered_output(4);
   bh4_w5_10 <= tile_10_filtered_output(5);
   bh4_w6_10 <= tile_10_filtered_output(6);
   bh4_w7_10 <= tile_10_filtered_output(7);
   bh4_w8_10 <= tile_10_filtered_output(8);
   bh4_w9_10 <= tile_10_filtered_output(9);
   bh4_w10_10 <= tile_10_filtered_output(10);
   bh4_w11_10 <= tile_10_filtered_output(11);
   bh4_w12_10 <= tile_10_filtered_output(12);
   bh4_w13_10 <= tile_10_filtered_output(13);
   tile_11_X <= X(9 downto 9);
   tile_11_Y <= Y(33 downto 20);
   tile_11_mult: DSPBlock_1x14_F125_uid28
      port map ( clk  => clk,
                 X => tile_11_X,
                 Y => tile_11_Y,
                 R => tile_11_output);

   tile_11_filtered_output <= unsigned(tile_11_output(13 downto 0));
   bh4_w0_11 <= tile_11_filtered_output(0);
   bh4_w1_11 <= tile_11_filtered_output(1);
   bh4_w2_11 <= tile_11_filtered_output(2);
   bh4_w3_11 <= tile_11_filtered_output(3);
   bh4_w4_11 <= tile_11_filtered_output(4);
   bh4_w5_11 <= tile_11_filtered_output(5);
   bh4_w6_11 <= tile_11_filtered_output(6);
   bh4_w7_11 <= tile_11_filtered_output(7);
   bh4_w8_11 <= tile_11_filtered_output(8);
   bh4_w9_11 <= tile_11_filtered_output(9);
   bh4_w10_11 <= tile_11_filtered_output(10);
   bh4_w11_11 <= tile_11_filtered_output(11);
   bh4_w12_11 <= tile_11_filtered_output(12);
   bh4_w13_11 <= tile_11_filtered_output(13);
   tile_12_X <= X(33 downto 21);
   tile_12_Y <= Y(8 downto 8);
   tile_12_mult: DSPBlock_13x1_F125_uid30
      port map ( clk  => clk,
                 X => tile_12_X,
                 Y => tile_12_Y,
                 R => tile_12_output);

   tile_12_filtered_output <= unsigned(tile_12_output(12 downto 0));
   bh4_w0_12 <= tile_12_filtered_output(0);
   bh4_w1_12 <= tile_12_filtered_output(1);
   bh4_w2_12 <= tile_12_filtered_output(2);
   bh4_w3_12 <= tile_12_filtered_output(3);
   bh4_w4_12 <= tile_12_filtered_output(4);
   bh4_w5_12 <= tile_12_filtered_output(5);
   bh4_w6_12 <= tile_12_filtered_output(6);
   bh4_w7_12 <= tile_12_filtered_output(7);
   bh4_w8_12 <= tile_12_filtered_output(8);
   bh4_w9_12 <= tile_12_filtered_output(9);
   bh4_w10_12 <= tile_12_filtered_output(10);
   bh4_w11_12 <= tile_12_filtered_output(11);
   bh4_w12_12 <= tile_12_filtered_output(12);
   tile_13_X <= X(8 downto 8);
   tile_13_Y <= Y(33 downto 21);
   tile_13_mult: DSPBlock_1x13_F125_uid32
      port map ( clk  => clk,
                 X => tile_13_X,
                 Y => tile_13_Y,
                 R => tile_13_output);

   tile_13_filtered_output <= unsigned(tile_13_output(12 downto 0));
   bh4_w0_13 <= tile_13_filtered_output(0);
   bh4_w1_13 <= tile_13_filtered_output(1);
   bh4_w2_13 <= tile_13_filtered_output(2);
   bh4_w3_13 <= tile_13_filtered_output(3);
   bh4_w4_13 <= tile_13_filtered_output(4);
   bh4_w5_13 <= tile_13_filtered_output(5);
   bh4_w6_13 <= tile_13_filtered_output(6);
   bh4_w7_13 <= tile_13_filtered_output(7);
   bh4_w8_13 <= tile_13_filtered_output(8);
   bh4_w9_13 <= tile_13_filtered_output(9);
   bh4_w10_13 <= tile_13_filtered_output(10);
   bh4_w11_13 <= tile_13_filtered_output(11);
   bh4_w12_13 <= tile_13_filtered_output(12);
   tile_14_X <= X(7 downto 7);
   tile_14_Y <= Y(33 downto 22);
   tile_14_mult: DSPBlock_1x12_F125_uid34
      port map ( clk  => clk,
                 X => tile_14_X,
                 Y => tile_14_Y,
                 R => tile_14_output);

   tile_14_filtered_output <= unsigned(tile_14_output(11 downto 0));
   bh4_w0_14 <= tile_14_filtered_output(0);
   bh4_w1_14 <= tile_14_filtered_output(1);
   bh4_w2_14 <= tile_14_filtered_output(2);
   bh4_w3_14 <= tile_14_filtered_output(3);
   bh4_w4_14 <= tile_14_filtered_output(4);
   bh4_w5_14 <= tile_14_filtered_output(5);
   bh4_w6_14 <= tile_14_filtered_output(6);
   bh4_w7_14 <= tile_14_filtered_output(7);
   bh4_w8_14 <= tile_14_filtered_output(8);
   bh4_w9_14 <= tile_14_filtered_output(9);
   bh4_w10_14 <= tile_14_filtered_output(10);
   bh4_w11_14 <= tile_14_filtered_output(11);
   tile_15_X <= X(33 downto 22);
   tile_15_Y <= Y(7 downto 7);
   tile_15_mult: DSPBlock_12x1_F125_uid36
      port map ( clk  => clk,
                 X => tile_15_X,
                 Y => tile_15_Y,
                 R => tile_15_output);

   tile_15_filtered_output <= unsigned(tile_15_output(11 downto 0));
   bh4_w0_15 <= tile_15_filtered_output(0);
   bh4_w1_15 <= tile_15_filtered_output(1);
   bh4_w2_15 <= tile_15_filtered_output(2);
   bh4_w3_15 <= tile_15_filtered_output(3);
   bh4_w4_15 <= tile_15_filtered_output(4);
   bh4_w5_15 <= tile_15_filtered_output(5);
   bh4_w6_15 <= tile_15_filtered_output(6);
   bh4_w7_15 <= tile_15_filtered_output(7);
   bh4_w8_15 <= tile_15_filtered_output(8);
   bh4_w9_15 <= tile_15_filtered_output(9);
   bh4_w10_15 <= tile_15_filtered_output(10);
   bh4_w11_15 <= tile_15_filtered_output(11);
   tile_16_X <= X(33 downto 23);
   tile_16_Y <= Y(6 downto 6);
   tile_16_mult: DSPBlock_11x1_F125_uid38
      port map ( clk  => clk,
                 X => tile_16_X,
                 Y => tile_16_Y,
                 R => tile_16_output);

   tile_16_filtered_output <= unsigned(tile_16_output(10 downto 0));
   bh4_w0_16 <= tile_16_filtered_output(0);
   bh4_w1_16 <= tile_16_filtered_output(1);
   bh4_w2_16 <= tile_16_filtered_output(2);
   bh4_w3_16 <= tile_16_filtered_output(3);
   bh4_w4_16 <= tile_16_filtered_output(4);
   bh4_w5_16 <= tile_16_filtered_output(5);
   bh4_w6_16 <= tile_16_filtered_output(6);
   bh4_w7_16 <= tile_16_filtered_output(7);
   bh4_w8_16 <= tile_16_filtered_output(8);
   bh4_w9_16 <= tile_16_filtered_output(9);
   bh4_w10_16 <= tile_16_filtered_output(10);
   tile_17_X <= X(6 downto 6);
   tile_17_Y <= Y(33 downto 23);
   tile_17_mult: DSPBlock_1x11_F125_uid40
      port map ( clk  => clk,
                 X => tile_17_X,
                 Y => tile_17_Y,
                 R => tile_17_output);

   tile_17_filtered_output <= unsigned(tile_17_output(10 downto 0));
   bh4_w0_17 <= tile_17_filtered_output(0);
   bh4_w1_17 <= tile_17_filtered_output(1);
   bh4_w2_17 <= tile_17_filtered_output(2);
   bh4_w3_17 <= tile_17_filtered_output(3);
   bh4_w4_17 <= tile_17_filtered_output(4);
   bh4_w5_17 <= tile_17_filtered_output(5);
   bh4_w6_17 <= tile_17_filtered_output(6);
   bh4_w7_17 <= tile_17_filtered_output(7);
   bh4_w8_17 <= tile_17_filtered_output(8);
   bh4_w9_17 <= tile_17_filtered_output(9);
   bh4_w10_17 <= tile_17_filtered_output(10);
   tile_18_X <= X(33 downto 24);
   tile_18_Y <= Y(5 downto 5);
   tile_18_mult: DSPBlock_10x1_F125_uid42
      port map ( clk  => clk,
                 X => tile_18_X,
                 Y => tile_18_Y,
                 R => tile_18_output);

   tile_18_filtered_output <= unsigned(tile_18_output(9 downto 0));
   bh4_w0_18 <= tile_18_filtered_output(0);
   bh4_w1_18 <= tile_18_filtered_output(1);
   bh4_w2_18 <= tile_18_filtered_output(2);
   bh4_w3_18 <= tile_18_filtered_output(3);
   bh4_w4_18 <= tile_18_filtered_output(4);
   bh4_w5_18 <= tile_18_filtered_output(5);
   bh4_w6_18 <= tile_18_filtered_output(6);
   bh4_w7_18 <= tile_18_filtered_output(7);
   bh4_w8_18 <= tile_18_filtered_output(8);
   bh4_w9_18 <= tile_18_filtered_output(9);
   tile_19_X <= X(5 downto 5);
   tile_19_Y <= Y(33 downto 24);
   tile_19_mult: DSPBlock_1x10_F125_uid44
      port map ( clk  => clk,
                 X => tile_19_X,
                 Y => tile_19_Y,
                 R => tile_19_output);

   tile_19_filtered_output <= unsigned(tile_19_output(9 downto 0));
   bh4_w0_19 <= tile_19_filtered_output(0);
   bh4_w1_19 <= tile_19_filtered_output(1);
   bh4_w2_19 <= tile_19_filtered_output(2);
   bh4_w3_19 <= tile_19_filtered_output(3);
   bh4_w4_19 <= tile_19_filtered_output(4);
   bh4_w5_19 <= tile_19_filtered_output(5);
   bh4_w6_19 <= tile_19_filtered_output(6);
   bh4_w7_19 <= tile_19_filtered_output(7);
   bh4_w8_19 <= tile_19_filtered_output(8);
   bh4_w9_19 <= tile_19_filtered_output(9);
   tile_20_X <= X(33 downto 25);
   tile_20_Y <= Y(4 downto 4);
   tile_20_mult: DSPBlock_9x1_F125_uid46
      port map ( clk  => clk,
                 X => tile_20_X,
                 Y => tile_20_Y,
                 R => tile_20_output);

   tile_20_filtered_output <= unsigned(tile_20_output(8 downto 0));
   bh4_w0_20 <= tile_20_filtered_output(0);
   bh4_w1_20 <= tile_20_filtered_output(1);
   bh4_w2_20 <= tile_20_filtered_output(2);
   bh4_w3_20 <= tile_20_filtered_output(3);
   bh4_w4_20 <= tile_20_filtered_output(4);
   bh4_w5_20 <= tile_20_filtered_output(5);
   bh4_w6_20 <= tile_20_filtered_output(6);
   bh4_w7_20 <= tile_20_filtered_output(7);
   bh4_w8_20 <= tile_20_filtered_output(8);
   tile_21_X <= X(4 downto 4);
   tile_21_Y <= Y(33 downto 25);
   tile_21_mult: DSPBlock_1x9_F125_uid48
      port map ( clk  => clk,
                 X => tile_21_X,
                 Y => tile_21_Y,
                 R => tile_21_output);

   tile_21_filtered_output <= unsigned(tile_21_output(8 downto 0));
   bh4_w0_21 <= tile_21_filtered_output(0);
   bh4_w1_21 <= tile_21_filtered_output(1);
   bh4_w2_21 <= tile_21_filtered_output(2);
   bh4_w3_21 <= tile_21_filtered_output(3);
   bh4_w4_21 <= tile_21_filtered_output(4);
   bh4_w5_21 <= tile_21_filtered_output(5);
   bh4_w6_21 <= tile_21_filtered_output(6);
   bh4_w7_21 <= tile_21_filtered_output(7);
   bh4_w8_21 <= tile_21_filtered_output(8);
   tile_22_X <= X(33 downto 26);
   tile_22_Y <= Y(3 downto 3);
   tile_22_mult: DSPBlock_8x1_F125_uid50
      port map ( clk  => clk,
                 X => tile_22_X,
                 Y => tile_22_Y,
                 R => tile_22_output);

   tile_22_filtered_output <= unsigned(tile_22_output(7 downto 0));
   bh4_w0_22 <= tile_22_filtered_output(0);
   bh4_w1_22 <= tile_22_filtered_output(1);
   bh4_w2_22 <= tile_22_filtered_output(2);
   bh4_w3_22 <= tile_22_filtered_output(3);
   bh4_w4_22 <= tile_22_filtered_output(4);
   bh4_w5_22 <= tile_22_filtered_output(5);
   bh4_w6_22 <= tile_22_filtered_output(6);
   bh4_w7_22 <= tile_22_filtered_output(7);
   tile_23_X <= X(3 downto 3);
   tile_23_Y <= Y(33 downto 26);
   tile_23_mult: DSPBlock_1x8_F125_uid52
      port map ( clk  => clk,
                 X => tile_23_X,
                 Y => tile_23_Y,
                 R => tile_23_output);

   tile_23_filtered_output <= unsigned(tile_23_output(7 downto 0));
   bh4_w0_23 <= tile_23_filtered_output(0);
   bh4_w1_23 <= tile_23_filtered_output(1);
   bh4_w2_23 <= tile_23_filtered_output(2);
   bh4_w3_23 <= tile_23_filtered_output(3);
   bh4_w4_23 <= tile_23_filtered_output(4);
   bh4_w5_23 <= tile_23_filtered_output(5);
   bh4_w6_23 <= tile_23_filtered_output(6);
   bh4_w7_23 <= tile_23_filtered_output(7);
   tile_24_X <= X(33 downto 27);
   tile_24_Y <= Y(2 downto 2);
   tile_24_mult: DSPBlock_7x1_F125_uid54
      port map ( clk  => clk,
                 X => tile_24_X,
                 Y => tile_24_Y,
                 R => tile_24_output);

   tile_24_filtered_output <= unsigned(tile_24_output(6 downto 0));
   bh4_w0_24 <= tile_24_filtered_output(0);
   bh4_w1_24 <= tile_24_filtered_output(1);
   bh4_w2_24 <= tile_24_filtered_output(2);
   bh4_w3_24 <= tile_24_filtered_output(3);
   bh4_w4_24 <= tile_24_filtered_output(4);
   bh4_w5_24 <= tile_24_filtered_output(5);
   bh4_w6_24 <= tile_24_filtered_output(6);
   tile_25_X <= X(2 downto 2);
   tile_25_Y <= Y(33 downto 27);
   tile_25_mult: DSPBlock_1x7_F125_uid56
      port map ( clk  => clk,
                 X => tile_25_X,
                 Y => tile_25_Y,
                 R => tile_25_output);

   tile_25_filtered_output <= unsigned(tile_25_output(6 downto 0));
   bh4_w0_25 <= tile_25_filtered_output(0);
   bh4_w1_25 <= tile_25_filtered_output(1);
   bh4_w2_25 <= tile_25_filtered_output(2);
   bh4_w3_25 <= tile_25_filtered_output(3);
   bh4_w4_25 <= tile_25_filtered_output(4);
   bh4_w5_25 <= tile_25_filtered_output(5);
   bh4_w6_25 <= tile_25_filtered_output(6);
   tile_26_X <= X(1 downto 1);
   tile_26_Y <= Y(33 downto 28);
   tile_26_mult: DSPBlock_1x6_F125_uid58
      port map ( clk  => clk,
                 X => tile_26_X,
                 Y => tile_26_Y,
                 R => tile_26_output);

   tile_26_filtered_output <= unsigned(tile_26_output(5 downto 0));
   bh4_w0_26 <= tile_26_filtered_output(0);
   bh4_w1_26 <= tile_26_filtered_output(1);
   bh4_w2_26 <= tile_26_filtered_output(2);
   bh4_w3_26 <= tile_26_filtered_output(3);
   bh4_w4_26 <= tile_26_filtered_output(4);
   bh4_w5_26 <= tile_26_filtered_output(5);
   tile_27_X <= X(0 downto 0);
   tile_27_Y <= Y(33 downto 29);
   tile_27_mult: DSPBlock_1x5_F125_uid60
      port map ( clk  => clk,
                 X => tile_27_X,
                 Y => tile_27_Y,
                 R => tile_27_output);

   tile_27_filtered_output <= unsigned(tile_27_output(4 downto 0));
   bh4_w0_27 <= tile_27_filtered_output(0);
   bh4_w1_27 <= tile_27_filtered_output(1);
   bh4_w2_27 <= tile_27_filtered_output(2);
   bh4_w3_27 <= tile_27_filtered_output(3);
   bh4_w4_27 <= tile_27_filtered_output(4);
   tile_28_X <= X(33 downto 29);
   tile_28_Y <= Y(1 downto 1);
   tile_28_mult: DSPBlock_5x1_F125_uid62
      port map ( clk  => clk,
                 X => tile_28_X,
                 Y => tile_28_Y,
                 R => tile_28_output);

   tile_28_filtered_output <= unsigned(tile_28_output(4 downto 0));
   bh4_w1_28 <= tile_28_filtered_output(0);
   bh4_w2_28 <= tile_28_filtered_output(1);
   bh4_w3_28 <= tile_28_filtered_output(2);
   bh4_w4_28 <= tile_28_filtered_output(3);
   bh4_w5_27 <= tile_28_filtered_output(4);
   tile_29_X <= X(33 downto 30);
   tile_29_Y <= Y(0 downto 0);
   tile_29_mult: DSPBlock_4x1_F125_uid64
      port map ( clk  => clk,
                 X => tile_29_X,
                 Y => tile_29_Y,
                 R => tile_29_output);

   tile_29_filtered_output <= unsigned(tile_29_output(3 downto 0));
   bh4_w1_29 <= tile_29_filtered_output(0);
   bh4_w2_29 <= tile_29_filtered_output(1);
   bh4_w3_29 <= tile_29_filtered_output(2);
   bh4_w4_29 <= tile_29_filtered_output(3);
   tile_30_X <= X(33 downto 31);
   tile_30_Y <= Y(33 downto 15);
   tile_30_mult: DSPBlock_3x19_F125_uid66
      port map ( clk  => clk,
                 X => tile_30_X,
                 Y => tile_30_Y,
                 R => tile_30_output);

   tile_30_filtered_output <= unsigned(tile_30_output(21 downto 0));
   bh4_w17_4 <= tile_30_filtered_output(0);
   bh4_w18_2 <= tile_30_filtered_output(1);
   bh4_w19_1 <= tile_30_filtered_output(2);
   bh4_w20_1 <= tile_30_filtered_output(3);
   bh4_w21_1 <= tile_30_filtered_output(4);
   bh4_w22_1 <= tile_30_filtered_output(5);
   bh4_w23_1 <= tile_30_filtered_output(6);
   bh4_w24_1 <= tile_30_filtered_output(7);
   bh4_w25_1 <= tile_30_filtered_output(8);
   bh4_w26_1 <= tile_30_filtered_output(9);
   bh4_w27_1 <= tile_30_filtered_output(10);
   bh4_w28_1 <= tile_30_filtered_output(11);
   bh4_w29_1 <= tile_30_filtered_output(12);
   bh4_w30_1 <= tile_30_filtered_output(13);
   bh4_w31_1 <= tile_30_filtered_output(14);
   bh4_w32_1 <= tile_30_filtered_output(15);
   bh4_w33_1 <= tile_30_filtered_output(16);
   bh4_w34_1 <= tile_30_filtered_output(17);
   bh4_w35_1 <= tile_30_filtered_output(18);
   bh4_w36_0 <= tile_30_filtered_output(19);
   bh4_w37_0 <= tile_30_filtered_output(20);
   bh4_w38_0 <= tile_30_filtered_output(21);

   -- Adding the constant bits
   bh4_w0_28 <= '1';
   bh4_w1_30 <= '1';
   bh4_w2_30 <= '1';
   bh4_w3_30 <= '1';
   bh4_w4_30 <= '1';


   Compressor_6_3_F125_uid69_bh4_uid70_In0 <= "" & bh4_w0_14 & bh4_w0_28 & bh4_w0_27 & bh4_w0_26 & bh4_w0_25 & bh4_w0_24;
   bh4_w0_29 <= Compressor_6_3_F125_uid69_bh4_uid70_Out0(0);
   bh4_w1_31 <= Compressor_6_3_F125_uid69_bh4_uid70_Out0(1);
   bh4_w2_31 <= Compressor_6_3_F125_uid69_bh4_uid70_Out0(2);
   Compressor_6_3_F125_uid69_uid70: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid70_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid70_Out0_copy71);
   Compressor_6_3_F125_uid69_bh4_uid70_Out0 <= Compressor_6_3_F125_uid69_bh4_uid70_Out0_copy71; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid72_In0 <= "" & bh4_w0_0 & bh4_w0_1 & bh4_w0_2 & bh4_w0_3 & bh4_w0_4 & bh4_w0_5;
   bh4_w0_30 <= Compressor_6_3_F125_uid69_bh4_uid72_Out0(0);
   bh4_w1_32 <= Compressor_6_3_F125_uid69_bh4_uid72_Out0(1);
   bh4_w2_32 <= Compressor_6_3_F125_uid69_bh4_uid72_Out0(2);
   Compressor_6_3_F125_uid69_uid72: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid72_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid72_Out0_copy73);
   Compressor_6_3_F125_uid69_bh4_uid72_Out0 <= Compressor_6_3_F125_uid69_bh4_uid72_Out0_copy73; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid74_In0 <= "" & bh4_w0_13 & bh4_w0_23 & bh4_w0_22 & bh4_w0_21 & bh4_w0_20 & bh4_w0_19;
   bh4_w0_31 <= Compressor_6_3_F125_uid69_bh4_uid74_Out0(0);
   bh4_w1_33 <= Compressor_6_3_F125_uid69_bh4_uid74_Out0(1);
   bh4_w2_33 <= Compressor_6_3_F125_uid69_bh4_uid74_Out0(2);
   Compressor_6_3_F125_uid69_uid74: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid74_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid74_Out0_copy75);
   Compressor_6_3_F125_uid69_bh4_uid74_Out0 <= Compressor_6_3_F125_uid69_bh4_uid74_Out0_copy75; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid76_In0 <= "" & bh4_w0_6 & bh4_w0_7 & bh4_w0_8 & bh4_w0_9 & bh4_w0_10 & bh4_w0_11;
   bh4_w0_32 <= Compressor_6_3_F125_uid69_bh4_uid76_Out0(0);
   bh4_w1_34 <= Compressor_6_3_F125_uid69_bh4_uid76_Out0(1);
   bh4_w2_34 <= Compressor_6_3_F125_uid69_bh4_uid76_Out0(2);
   Compressor_6_3_F125_uid69_uid76: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid76_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid76_Out0_copy77);
   Compressor_6_3_F125_uid69_bh4_uid76_Out0 <= Compressor_6_3_F125_uid69_bh4_uid76_Out0_copy77; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid80_In0 <= "" & bh4_w0_15 & bh4_w0_16 & bh4_w0_17 & bh4_w0_18;
   Compressor_14_3_F125_uid79_bh4_uid80_In1 <= "" & bh4_w1_22;
   bh4_w0_33 <= Compressor_14_3_F125_uid79_bh4_uid80_Out0(0);
   bh4_w1_35 <= Compressor_14_3_F125_uid79_bh4_uid80_Out0(1);
   bh4_w2_35 <= Compressor_14_3_F125_uid79_bh4_uid80_Out0(2);
   Compressor_14_3_F125_uid79_uid80: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid80_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid80_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid80_Out0_copy81);
   Compressor_14_3_F125_uid79_bh4_uid80_Out0 <= Compressor_14_3_F125_uid79_bh4_uid80_Out0_copy81; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid82_In0 <= "" & bh4_w1_6 & bh4_w1_0 & bh4_w1_13 & bh4_w1_12 & bh4_w1_11 & bh4_w1_10;
   bh4_w1_36 <= Compressor_6_3_F125_uid69_bh4_uid82_Out0(0);
   bh4_w2_36 <= Compressor_6_3_F125_uid69_bh4_uid82_Out0(1);
   bh4_w3_31 <= Compressor_6_3_F125_uid69_bh4_uid82_Out0(2);
   Compressor_6_3_F125_uid69_uid82: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid82_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid82_Out0_copy83);
   Compressor_6_3_F125_uid69_bh4_uid82_Out0 <= Compressor_6_3_F125_uid69_bh4_uid82_Out0_copy83; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid84_In0 <= "" & bh4_w1_14 & bh4_w1_15 & bh4_w1_16 & bh4_w1_17 & bh4_w1_18 & bh4_w1_19;
   bh4_w1_37 <= Compressor_6_3_F125_uid69_bh4_uid84_Out0(0);
   bh4_w2_37 <= Compressor_6_3_F125_uid69_bh4_uid84_Out0(1);
   bh4_w3_32 <= Compressor_6_3_F125_uid69_bh4_uid84_Out0(2);
   Compressor_6_3_F125_uid69_uid84: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid84_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid84_Out0_copy85);
   Compressor_6_3_F125_uid69_bh4_uid84_Out0 <= Compressor_6_3_F125_uid69_bh4_uid84_Out0_copy85; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid86_In0 <= "" & bh4_w1_30 & bh4_w1_9 & bh4_w1_8 & bh4_w1_7 & bh4_w1_29 & bh4_w1_5;
   bh4_w1_38 <= Compressor_6_3_F125_uid69_bh4_uid86_Out0(0);
   bh4_w2_38 <= Compressor_6_3_F125_uid69_bh4_uid86_Out0(1);
   bh4_w3_33 <= Compressor_6_3_F125_uid69_bh4_uid86_Out0(2);
   Compressor_6_3_F125_uid69_uid86: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid86_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid86_Out0_copy87);
   Compressor_6_3_F125_uid69_bh4_uid86_Out0 <= Compressor_6_3_F125_uid69_bh4_uid86_Out0_copy87; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid88_In0 <= "" & bh4_w1_20 & bh4_w1_21 & bh4_w1_23 & bh4_w1_24 & bh4_w1_25 & bh4_w1_26;
   bh4_w1_39 <= Compressor_6_3_F125_uid69_bh4_uid88_Out0(0);
   bh4_w2_39 <= Compressor_6_3_F125_uid69_bh4_uid88_Out0(1);
   bh4_w3_34 <= Compressor_6_3_F125_uid69_bh4_uid88_Out0(2);
   Compressor_6_3_F125_uid69_uid88: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid88_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid88_Out0_copy89);
   Compressor_6_3_F125_uid69_bh4_uid88_Out0 <= Compressor_6_3_F125_uid69_bh4_uid88_Out0_copy89; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid90_In0 <= "" & bh4_w1_28 & bh4_w1_4 & bh4_w1_3 & bh4_w1_2 & bh4_w1_1 & bh4_w1_27;
   bh4_w1_40 <= Compressor_6_3_F125_uid69_bh4_uid90_Out0(0);
   bh4_w2_40 <= Compressor_6_3_F125_uid69_bh4_uid90_Out0(1);
   bh4_w3_35 <= Compressor_6_3_F125_uid69_bh4_uid90_Out0(2);
   Compressor_6_3_F125_uid69_uid90: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid90_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid90_Out0_copy91);
   Compressor_6_3_F125_uid69_bh4_uid90_Out0 <= Compressor_6_3_F125_uid69_bh4_uid90_Out0_copy91; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid92_In0 <= "" & bh4_w2_20 & bh4_w2_19 & bh4_w2_21 & bh4_w2_14 & bh4_w2_15 & bh4_w2_16;
   bh4_w2_41 <= Compressor_6_3_F125_uid69_bh4_uid92_Out0(0);
   bh4_w3_36 <= Compressor_6_3_F125_uid69_bh4_uid92_Out0(1);
   bh4_w4_31 <= Compressor_6_3_F125_uid69_bh4_uid92_Out0(2);
   Compressor_6_3_F125_uid69_uid92: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid92_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid92_Out0_copy93);
   Compressor_6_3_F125_uid69_bh4_uid92_Out0 <= Compressor_6_3_F125_uid69_bh4_uid92_Out0_copy93; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid94_In0 <= "" & bh4_w2_7 & bh4_w2_28 & bh4_w2_29 & bh4_w2_30 & bh4_w2_0 & bh4_w2_13;
   bh4_w2_42 <= Compressor_6_3_F125_uid69_bh4_uid94_Out0(0);
   bh4_w3_37 <= Compressor_6_3_F125_uid69_bh4_uid94_Out0(1);
   bh4_w4_32 <= Compressor_6_3_F125_uid69_bh4_uid94_Out0(2);
   Compressor_6_3_F125_uid69_uid94: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid94_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid94_Out0_copy95);
   Compressor_6_3_F125_uid69_bh4_uid94_Out0 <= Compressor_6_3_F125_uid69_bh4_uid94_Out0_copy95; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid96_In0 <= "" & bh4_w2_17 & bh4_w2_18 & bh4_w2_22 & bh4_w2_23 & bh4_w2_24 & bh4_w2_25;
   bh4_w2_43 <= Compressor_6_3_F125_uid69_bh4_uid96_Out0(0);
   bh4_w3_38 <= Compressor_6_3_F125_uid69_bh4_uid96_Out0(1);
   bh4_w4_33 <= Compressor_6_3_F125_uid69_bh4_uid96_Out0(2);
   Compressor_6_3_F125_uid69_uid96: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid96_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid96_Out0_copy97);
   Compressor_6_3_F125_uid69_bh4_uid96_Out0 <= Compressor_6_3_F125_uid69_bh4_uid96_Out0_copy97; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid98_In0 <= "" & bh4_w2_8 & bh4_w2_27 & bh4_w2_12 & bh4_w2_11 & bh4_w2_10 & bh4_w2_9;
   bh4_w2_44 <= Compressor_6_3_F125_uid69_bh4_uid98_Out0(0);
   bh4_w3_39 <= Compressor_6_3_F125_uid69_bh4_uid98_Out0(1);
   bh4_w4_34 <= Compressor_6_3_F125_uid69_bh4_uid98_Out0(2);
   Compressor_6_3_F125_uid69_uid98: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid98_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid98_Out0_copy99);
   Compressor_6_3_F125_uid69_bh4_uid98_Out0 <= Compressor_6_3_F125_uid69_bh4_uid98_Out0_copy99; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid100_In0 <= "" & bh4_w2_26 & bh4_w2_6 & bh4_w2_5 & bh4_w2_4 & bh4_w2_3 & bh4_w2_2;
   bh4_w2_45 <= Compressor_6_3_F125_uid69_bh4_uid100_Out0(0);
   bh4_w3_40 <= Compressor_6_3_F125_uid69_bh4_uid100_Out0(1);
   bh4_w4_35 <= Compressor_6_3_F125_uid69_bh4_uid100_Out0(2);
   Compressor_6_3_F125_uid69_uid100: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid100_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid100_Out0_copy101);
   Compressor_6_3_F125_uid69_bh4_uid100_Out0 <= Compressor_6_3_F125_uid69_bh4_uid100_Out0_copy101; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid102_In0 <= "" & bh4_w3_11 & bh4_w3_12 & bh4_w3_10 & bh4_w3_17 & bh4_w3_0 & bh4_w3_15;
   bh4_w3_41 <= Compressor_6_3_F125_uid69_bh4_uid102_Out0(0);
   bh4_w4_36 <= Compressor_6_3_F125_uid69_bh4_uid102_Out0(1);
   bh4_w5_28 <= Compressor_6_3_F125_uid69_bh4_uid102_Out0(2);
   Compressor_6_3_F125_uid69_uid102: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid102_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid102_Out0_copy103);
   Compressor_6_3_F125_uid69_bh4_uid102_Out0 <= Compressor_6_3_F125_uid69_bh4_uid102_Out0_copy103; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid104_In0 <= "" & bh4_w3_24 & bh4_w3_3 & bh4_w3_2 & bh4_w3_1 & bh4_w3_16 & bh4_w3_18;
   bh4_w3_42 <= Compressor_6_3_F125_uid69_bh4_uid104_Out0(0);
   bh4_w4_37 <= Compressor_6_3_F125_uid69_bh4_uid104_Out0(1);
   bh4_w5_29 <= Compressor_6_3_F125_uid69_bh4_uid104_Out0(2);
   Compressor_6_3_F125_uid69_uid104: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid104_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid104_Out0_copy105);
   Compressor_6_3_F125_uid69_bh4_uid104_Out0 <= Compressor_6_3_F125_uid69_bh4_uid104_Out0_copy105; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid106_In0 <= "" & bh4_w3_14 & bh4_w3_13 & bh4_w3_9 & bh4_w3_8 & bh4_w3_7 & bh4_w3_6;
   bh4_w3_43 <= Compressor_6_3_F125_uid69_bh4_uid106_Out0(0);
   bh4_w4_38 <= Compressor_6_3_F125_uid69_bh4_uid106_Out0(1);
   bh4_w5_30 <= Compressor_6_3_F125_uid69_bh4_uid106_Out0(2);
   Compressor_6_3_F125_uid69_uid106: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid106_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid106_Out0_copy107);
   Compressor_6_3_F125_uid69_bh4_uid106_Out0 <= Compressor_6_3_F125_uid69_bh4_uid106_Out0_copy107; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid108_In0 <= "" & bh4_w3_23 & bh4_w3_4 & bh4_w3_19 & bh4_w3_20 & bh4_w3_21 & bh4_w3_22;
   bh4_w3_44 <= Compressor_6_3_F125_uid69_bh4_uid108_Out0(0);
   bh4_w4_39 <= Compressor_6_3_F125_uid69_bh4_uid108_Out0(1);
   bh4_w5_31 <= Compressor_6_3_F125_uid69_bh4_uid108_Out0(2);
   Compressor_6_3_F125_uid69_uid108: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid108_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid108_Out0_copy109);
   Compressor_6_3_F125_uid69_bh4_uid108_Out0 <= Compressor_6_3_F125_uid69_bh4_uid108_Out0_copy109; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid110_In0 <= "" & bh4_w3_5 & bh4_w3_25 & bh4_w3_26 & bh4_w3_27 & bh4_w3_28 & bh4_w3_29;
   bh4_w3_45 <= Compressor_6_3_F125_uid69_bh4_uid110_Out0(0);
   bh4_w4_40 <= Compressor_6_3_F125_uid69_bh4_uid110_Out0(1);
   bh4_w5_32 <= Compressor_6_3_F125_uid69_bh4_uid110_Out0(2);
   Compressor_6_3_F125_uid69_uid110: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid110_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid110_Out0_copy111);
   Compressor_6_3_F125_uid69_bh4_uid110_Out0 <= Compressor_6_3_F125_uid69_bh4_uid110_Out0_copy111; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid112_In0 <= "" & bh4_w4_20 & bh4_w4_19 & bh4_w4_21 & bh4_w4_14 & bh4_w4_16 & bh4_w4_0;
   bh4_w4_41 <= Compressor_6_3_F125_uid69_bh4_uid112_Out0(0);
   bh4_w5_33 <= Compressor_6_3_F125_uid69_bh4_uid112_Out0(1);
   bh4_w6_26 <= Compressor_6_3_F125_uid69_bh4_uid112_Out0(2);
   Compressor_6_3_F125_uid69_uid112: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid112_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid112_Out0_copy113);
   Compressor_6_3_F125_uid69_bh4_uid112_Out0 <= Compressor_6_3_F125_uid69_bh4_uid112_Out0_copy113; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid114_In0 <= "" & bh4_w4_7 & bh4_w4_28 & bh4_w4_29 & bh4_w4_30 & bh4_w4_15 & bh4_w4_13;
   bh4_w4_42 <= Compressor_6_3_F125_uid69_bh4_uid114_Out0(0);
   bh4_w5_34 <= Compressor_6_3_F125_uid69_bh4_uid114_Out0(1);
   bh4_w6_27 <= Compressor_6_3_F125_uid69_bh4_uid114_Out0(2);
   Compressor_6_3_F125_uid69_uid114: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid114_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid114_Out0_copy115);
   Compressor_6_3_F125_uid69_bh4_uid114_Out0 <= Compressor_6_3_F125_uid69_bh4_uid114_Out0_copy115; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid116_In0 <= "" & bh4_w4_17 & bh4_w4_18 & bh4_w4_22 & bh4_w4_23 & bh4_w4_24 & bh4_w4_25;
   bh4_w4_43 <= Compressor_6_3_F125_uid69_bh4_uid116_Out0(0);
   bh4_w5_35 <= Compressor_6_3_F125_uid69_bh4_uid116_Out0(1);
   bh4_w6_28 <= Compressor_6_3_F125_uid69_bh4_uid116_Out0(2);
   Compressor_6_3_F125_uid69_uid116: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid116_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid116_Out0_copy117);
   Compressor_6_3_F125_uid69_bh4_uid116_Out0 <= Compressor_6_3_F125_uid69_bh4_uid116_Out0_copy117; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid118_In0 <= "" & bh4_w4_8 & bh4_w4_27 & bh4_w4_12 & bh4_w4_11 & bh4_w4_10 & bh4_w4_9;
   bh4_w4_44 <= Compressor_6_3_F125_uid69_bh4_uid118_Out0(0);
   bh4_w5_36 <= Compressor_6_3_F125_uid69_bh4_uid118_Out0(1);
   bh4_w6_29 <= Compressor_6_3_F125_uid69_bh4_uid118_Out0(2);
   Compressor_6_3_F125_uid69_uid118: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid118_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid118_Out0_copy119);
   Compressor_6_3_F125_uid69_bh4_uid118_Out0 <= Compressor_6_3_F125_uid69_bh4_uid118_Out0_copy119; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid120_In0 <= "" & bh4_w4_26 & bh4_w4_6 & bh4_w4_5 & bh4_w4_4 & bh4_w4_3 & bh4_w4_2;
   bh4_w4_45 <= Compressor_6_3_F125_uid69_bh4_uid120_Out0(0);
   bh4_w5_37 <= Compressor_6_3_F125_uid69_bh4_uid120_Out0(1);
   bh4_w6_30 <= Compressor_6_3_F125_uid69_bh4_uid120_Out0(2);
   Compressor_6_3_F125_uid69_uid120: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid120_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid120_Out0_copy121);
   Compressor_6_3_F125_uid69_bh4_uid120_Out0 <= Compressor_6_3_F125_uid69_bh4_uid120_Out0_copy121; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid122_In0 <= "" & bh4_w5_9 & bh4_w5_10 & bh4_w5_16 & bh4_w5_15 & bh4_w5_0 & bh4_w5_13;
   bh4_w5_38 <= Compressor_6_3_F125_uid69_bh4_uid122_Out0(0);
   bh4_w6_31 <= Compressor_6_3_F125_uid69_bh4_uid122_Out0(1);
   bh4_w7_24 <= Compressor_6_3_F125_uid69_bh4_uid122_Out0(2);
   Compressor_6_3_F125_uid69_uid122: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid122_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid122_Out0_copy123);
   Compressor_6_3_F125_uid69_bh4_uid122_Out0 <= Compressor_6_3_F125_uid69_bh4_uid122_Out0_copy123; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid124_In0 <= "" & bh4_w5_23 & bh4_w5_2 & bh4_w5_1 & bh4_w5_14 & bh4_w5_17 & bh4_w5_18;
   bh4_w5_39 <= Compressor_6_3_F125_uid69_bh4_uid124_Out0(0);
   bh4_w6_32 <= Compressor_6_3_F125_uid69_bh4_uid124_Out0(1);
   bh4_w7_25 <= Compressor_6_3_F125_uid69_bh4_uid124_Out0(2);
   Compressor_6_3_F125_uid69_uid124: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid124_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid124_Out0_copy125);
   Compressor_6_3_F125_uid69_bh4_uid124_Out0 <= Compressor_6_3_F125_uid69_bh4_uid124_Out0_copy125; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid126_In0 <= "" & bh4_w5_12 & bh4_w5_11 & bh4_w5_8 & bh4_w5_7 & bh4_w5_6 & bh4_w5_5;
   bh4_w5_40 <= Compressor_6_3_F125_uid69_bh4_uid126_Out0(0);
   bh4_w6_33 <= Compressor_6_3_F125_uid69_bh4_uid126_Out0(1);
   bh4_w7_26 <= Compressor_6_3_F125_uid69_bh4_uid126_Out0(2);
   Compressor_6_3_F125_uid69_uid126: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid126_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid126_Out0_copy127);
   Compressor_6_3_F125_uid69_bh4_uid126_Out0 <= Compressor_6_3_F125_uid69_bh4_uid126_Out0_copy127; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid128_In0 <= "" & bh4_w5_3 & bh4_w5_19 & bh4_w5_20 & bh4_w5_21 & bh4_w5_22 & bh4_w5_4;
   bh4_w5_41 <= Compressor_6_3_F125_uid69_bh4_uid128_Out0(0);
   bh4_w6_34 <= Compressor_6_3_F125_uid69_bh4_uid128_Out0(1);
   bh4_w7_27 <= Compressor_6_3_F125_uid69_bh4_uid128_Out0(2);
   Compressor_6_3_F125_uid69_uid128: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid128_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid128_Out0_copy129);
   Compressor_6_3_F125_uid69_bh4_uid128_Out0 <= Compressor_6_3_F125_uid69_bh4_uid128_Out0_copy129; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid130_In0 <= "" & bh4_w5_24 & bh4_w5_25 & bh4_w5_26 & bh4_w5_27;
   Compressor_14_3_F125_uid79_bh4_uid130_In1 <= "" & bh4_w6_2;
   bh4_w5_42 <= Compressor_14_3_F125_uid79_bh4_uid130_Out0(0);
   bh4_w6_35 <= Compressor_14_3_F125_uid79_bh4_uid130_Out0(1);
   bh4_w7_28 <= Compressor_14_3_F125_uid79_bh4_uid130_Out0(2);
   Compressor_14_3_F125_uid79_uid130: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid130_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid130_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid130_Out0_copy131);
   Compressor_14_3_F125_uid79_bh4_uid130_Out0 <= Compressor_14_3_F125_uid79_bh4_uid130_Out0_copy131; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid132_In0 <= "" & bh4_w6_17 & bh4_w6_10 & bh4_w6_11 & bh4_w6_12 & bh4_w6_13 & bh4_w6_14;
   bh4_w6_36 <= Compressor_6_3_F125_uid69_bh4_uid132_Out0(0);
   bh4_w7_29 <= Compressor_6_3_F125_uid69_bh4_uid132_Out0(1);
   bh4_w8_22 <= Compressor_6_3_F125_uid69_bh4_uid132_Out0(2);
   Compressor_6_3_F125_uid69_uid132: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid132_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid132_Out0_copy133);
   Compressor_6_3_F125_uid69_bh4_uid132_Out0 <= Compressor_6_3_F125_uid69_bh4_uid132_Out0_copy133; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid134_In0 <= "" & bh4_w6_25 & bh4_w6_0 & bh4_w6_9 & bh4_w6_8 & bh4_w6_7 & bh4_w6_6;
   bh4_w6_37 <= Compressor_6_3_F125_uid69_bh4_uid134_Out0(0);
   bh4_w7_30 <= Compressor_6_3_F125_uid69_bh4_uid134_Out0(1);
   bh4_w8_23 <= Compressor_6_3_F125_uid69_bh4_uid134_Out0(2);
   Compressor_6_3_F125_uid69_uid134: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid134_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid134_Out0_copy135);
   Compressor_6_3_F125_uid69_bh4_uid134_Out0 <= Compressor_6_3_F125_uid69_bh4_uid134_Out0_copy135; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid136_In0 <= "" & bh4_w6_16 & bh4_w6_15 & bh4_w6_18 & bh4_w6_19 & bh4_w6_20 & bh4_w6_21;
   bh4_w6_38 <= Compressor_6_3_F125_uid69_bh4_uid136_Out0(0);
   bh4_w7_31 <= Compressor_6_3_F125_uid69_bh4_uid136_Out0(1);
   bh4_w8_24 <= Compressor_6_3_F125_uid69_bh4_uid136_Out0(2);
   Compressor_6_3_F125_uid69_uid136: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid136_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid136_Out0_copy137);
   Compressor_6_3_F125_uid69_bh4_uid136_Out0 <= Compressor_6_3_F125_uid69_bh4_uid136_Out0_copy137; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid138_In0 <= "" & bh4_w6_3 & bh4_w6_24 & bh4_w6_5 & bh4_w6_4 & bh4_w6_23 & bh4_w6_1;
   bh4_w6_39 <= Compressor_6_3_F125_uid69_bh4_uid138_Out0(0);
   bh4_w7_32 <= Compressor_6_3_F125_uid69_bh4_uid138_Out0(1);
   bh4_w8_25 <= Compressor_6_3_F125_uid69_bh4_uid138_Out0(2);
   Compressor_6_3_F125_uid69_uid138: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid138_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid138_Out0_copy139);
   Compressor_6_3_F125_uid69_bh4_uid138_Out0 <= Compressor_6_3_F125_uid69_bh4_uid138_Out0_copy139; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid140_In0 <= "" & bh4_w7_17 & bh4_w7_18 & bh4_w7_19 & bh4_w7_20 & bh4_w7_21 & bh4_w7_22;
   bh4_w7_33 <= Compressor_6_3_F125_uid69_bh4_uid140_Out0(0);
   bh4_w8_26 <= Compressor_6_3_F125_uid69_bh4_uid140_Out0(1);
   bh4_w9_20 <= Compressor_6_3_F125_uid69_bh4_uid140_Out0(2);
   Compressor_6_3_F125_uid69_uid140: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid140_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid140_Out0_copy141);
   Compressor_6_3_F125_uid69_bh4_uid140_Out0 <= Compressor_6_3_F125_uid69_bh4_uid140_Out0_copy141; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid142_In0 <= "" & bh4_w7_8 & bh4_w7_16 & bh4_w7_15 & bh4_w7_14 & bh4_w7_13 & bh4_w7_0;
   bh4_w7_34 <= Compressor_6_3_F125_uid69_bh4_uid142_Out0(0);
   bh4_w8_27 <= Compressor_6_3_F125_uid69_bh4_uid142_Out0(1);
   bh4_w9_21 <= Compressor_6_3_F125_uid69_bh4_uid142_Out0(2);
   Compressor_6_3_F125_uid69_uid142: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid142_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid142_Out0_copy143);
   Compressor_6_3_F125_uid69_bh4_uid142_Out0 <= Compressor_6_3_F125_uid69_bh4_uid142_Out0_copy143; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid144_In0 <= "" & bh4_w7_23 & bh4_w7_1 & bh4_w7_12 & bh4_w7_11 & bh4_w7_10 & bh4_w7_9;
   bh4_w7_35 <= Compressor_6_3_F125_uid69_bh4_uid144_Out0(0);
   bh4_w8_28 <= Compressor_6_3_F125_uid69_bh4_uid144_Out0(1);
   bh4_w9_22 <= Compressor_6_3_F125_uid69_bh4_uid144_Out0(2);
   Compressor_6_3_F125_uid69_uid144: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid144_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid144_Out0_copy145);
   Compressor_6_3_F125_uid69_bh4_uid144_Out0 <= Compressor_6_3_F125_uid69_bh4_uid144_Out0_copy145; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid146_In0 <= "" & bh4_w7_7 & bh4_w7_6 & bh4_w7_5 & bh4_w7_4 & bh4_w7_3 & bh4_w7_2;
   bh4_w7_36 <= Compressor_6_3_F125_uid69_bh4_uid146_Out0(0);
   bh4_w8_29 <= Compressor_6_3_F125_uid69_bh4_uid146_Out0(1);
   bh4_w9_23 <= Compressor_6_3_F125_uid69_bh4_uid146_Out0(2);
   Compressor_6_3_F125_uid69_uid146: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid146_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid146_Out0_copy147);
   Compressor_6_3_F125_uid69_bh4_uid146_Out0 <= Compressor_6_3_F125_uid69_bh4_uid146_Out0_copy147; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid148_In0 <= "" & bh4_w8_7 & bh4_w8_21 & bh4_w8_20 & bh4_w8_19 & bh4_w8_18 & bh4_w8_17;
   bh4_w8_30 <= Compressor_6_3_F125_uid69_bh4_uid148_Out0(0);
   bh4_w9_24 <= Compressor_6_3_F125_uid69_bh4_uid148_Out0(1);
   bh4_w10_18 <= Compressor_6_3_F125_uid69_bh4_uid148_Out0(2);
   Compressor_6_3_F125_uid69_uid148: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid148_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid148_Out0_copy149);
   Compressor_6_3_F125_uid69_bh4_uid148_Out0 <= Compressor_6_3_F125_uid69_bh4_uid148_Out0_copy149; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid150_In0 <= "" & bh4_w8_0 & bh4_w8_1 & bh4_w8_2 & bh4_w8_3 & bh4_w8_4 & bh4_w8_5;
   bh4_w8_31 <= Compressor_6_3_F125_uid69_bh4_uid150_Out0(0);
   bh4_w9_25 <= Compressor_6_3_F125_uid69_bh4_uid150_Out0(1);
   bh4_w10_19 <= Compressor_6_3_F125_uid69_bh4_uid150_Out0(2);
   Compressor_6_3_F125_uid69_uid150: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid150_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid150_Out0_copy151);
   Compressor_6_3_F125_uid69_bh4_uid150_Out0 <= Compressor_6_3_F125_uid69_bh4_uid150_Out0_copy151; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid152_In0 <= "" & bh4_w8_6 & bh4_w8_16 & bh4_w8_15 & bh4_w8_14 & bh4_w8_13 & bh4_w8_12;
   bh4_w8_32 <= Compressor_6_3_F125_uid69_bh4_uid152_Out0(0);
   bh4_w9_26 <= Compressor_6_3_F125_uid69_bh4_uid152_Out0(1);
   bh4_w10_20 <= Compressor_6_3_F125_uid69_bh4_uid152_Out0(2);
   Compressor_6_3_F125_uid69_uid152: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid152_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid152_Out0_copy153);
   Compressor_6_3_F125_uid69_bh4_uid152_Out0 <= Compressor_6_3_F125_uid69_bh4_uid152_Out0_copy153; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid154_In0 <= "" & bh4_w8_8 & bh4_w8_9 & bh4_w8_10 & bh4_w8_11;
   Compressor_14_3_F125_uid79_bh4_uid154_In1 <= "" & bh4_w9_0;
   bh4_w8_33 <= Compressor_14_3_F125_uid79_bh4_uid154_Out0(0);
   bh4_w9_27 <= Compressor_14_3_F125_uid79_bh4_uid154_Out0(1);
   bh4_w10_21 <= Compressor_14_3_F125_uid79_bh4_uid154_Out0(2);
   Compressor_14_3_F125_uid79_uid154: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid154_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid154_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid154_Out0_copy155);
   Compressor_14_3_F125_uid79_bh4_uid154_Out0 <= Compressor_14_3_F125_uid79_bh4_uid154_Out0_copy155; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid156_In0 <= "" & bh4_w9_6 & bh4_w9_19 & bh4_w9_18 & bh4_w9_17 & bh4_w9_16 & bh4_w9_15;
   bh4_w9_28 <= Compressor_6_3_F125_uid69_bh4_uid156_Out0(0);
   bh4_w10_22 <= Compressor_6_3_F125_uid69_bh4_uid156_Out0(1);
   bh4_w11_16 <= Compressor_6_3_F125_uid69_bh4_uid156_Out0(2);
   Compressor_6_3_F125_uid69_uid156: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid156_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid156_Out0_copy157);
   Compressor_6_3_F125_uid69_bh4_uid156_Out0 <= Compressor_6_3_F125_uid69_bh4_uid156_Out0_copy157; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid158_In0 <= "" & bh4_w9_1 & bh4_w9_2 & bh4_w9_3 & bh4_w9_4 & bh4_w9_5 & bh4_w9_7;
   bh4_w9_29 <= Compressor_6_3_F125_uid69_bh4_uid158_Out0(0);
   bh4_w10_23 <= Compressor_6_3_F125_uid69_bh4_uid158_Out0(1);
   bh4_w11_17 <= Compressor_6_3_F125_uid69_bh4_uid158_Out0(2);
   Compressor_6_3_F125_uid69_uid158: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid158_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid158_Out0_copy159);
   Compressor_6_3_F125_uid69_bh4_uid158_Out0 <= Compressor_6_3_F125_uid69_bh4_uid158_Out0_copy159; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid160_In0 <= "" & bh4_w9_14 & bh4_w9_13 & bh4_w9_12 & bh4_w9_11 & bh4_w9_10 & bh4_w9_9;
   bh4_w9_30 <= Compressor_6_3_F125_uid69_bh4_uid160_Out0(0);
   bh4_w10_24 <= Compressor_6_3_F125_uid69_bh4_uid160_Out0(1);
   bh4_w11_18 <= Compressor_6_3_F125_uid69_bh4_uid160_Out0(2);
   Compressor_6_3_F125_uid69_uid160: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid160_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid160_Out0_copy161);
   Compressor_6_3_F125_uid69_bh4_uid160_Out0 <= Compressor_6_3_F125_uid69_bh4_uid160_Out0_copy161; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid162_In0 <= "" & bh4_w10_0 & bh4_w10_1 & bh4_w10_2 & bh4_w10_3 & bh4_w10_4 & bh4_w10_5;
   bh4_w10_25 <= Compressor_6_3_F125_uid69_bh4_uid162_Out0(0);
   bh4_w11_19 <= Compressor_6_3_F125_uid69_bh4_uid162_Out0(1);
   bh4_w12_14 <= Compressor_6_3_F125_uid69_bh4_uid162_Out0(2);
   Compressor_6_3_F125_uid69_uid162: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid162_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid162_Out0_copy163);
   Compressor_6_3_F125_uid69_bh4_uid162_Out0 <= Compressor_6_3_F125_uid69_bh4_uid162_Out0_copy163; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid164_In0 <= "" & bh4_w10_17 & bh4_w10_16 & bh4_w10_15 & bh4_w10_14 & bh4_w10_13 & bh4_w10_12;
   bh4_w10_26 <= Compressor_6_3_F125_uid69_bh4_uid164_Out0(0);
   bh4_w11_20 <= Compressor_6_3_F125_uid69_bh4_uid164_Out0(1);
   bh4_w12_15 <= Compressor_6_3_F125_uid69_bh4_uid164_Out0(2);
   Compressor_6_3_F125_uid69_uid164: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid164_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid164_Out0_copy165);
   Compressor_6_3_F125_uid69_bh4_uid164_Out0 <= Compressor_6_3_F125_uid69_bh4_uid164_Out0_copy165; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid166_In0 <= "" & bh4_w10_6 & bh4_w10_7 & bh4_w10_8 & bh4_w10_9 & bh4_w10_10 & bh4_w10_11;
   bh4_w10_27 <= Compressor_6_3_F125_uid69_bh4_uid166_Out0(0);
   bh4_w11_21 <= Compressor_6_3_F125_uid69_bh4_uid166_Out0(1);
   bh4_w12_16 <= Compressor_6_3_F125_uid69_bh4_uid166_Out0(2);
   Compressor_6_3_F125_uid69_uid166: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid166_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid166_Out0_copy167);
   Compressor_6_3_F125_uid69_bh4_uid166_Out0 <= Compressor_6_3_F125_uid69_bh4_uid166_Out0_copy167; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid168_In0 <= "" & bh4_w11_11 & bh4_w11_1 & bh4_w11_2 & bh4_w11_3 & bh4_w11_4 & bh4_w11_5;
   bh4_w11_22 <= Compressor_6_3_F125_uid69_bh4_uid168_Out0(0);
   bh4_w12_17 <= Compressor_6_3_F125_uid69_bh4_uid168_Out0(1);
   bh4_w13_12 <= Compressor_6_3_F125_uid69_bh4_uid168_Out0(2);
   Compressor_6_3_F125_uid69_uid168: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid168_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid168_Out0_copy169);
   Compressor_6_3_F125_uid69_bh4_uid168_Out0 <= Compressor_6_3_F125_uid69_bh4_uid168_Out0_copy169; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid170_In0 <= "" & bh4_w11_8 & bh4_w11_15 & bh4_w11_14 & bh4_w11_13 & bh4_w11_12 & bh4_w11_10;
   bh4_w11_23 <= Compressor_6_3_F125_uid69_bh4_uid170_Out0(0);
   bh4_w12_18 <= Compressor_6_3_F125_uid69_bh4_uid170_Out0(1);
   bh4_w13_13 <= Compressor_6_3_F125_uid69_bh4_uid170_Out0(2);
   Compressor_6_3_F125_uid69_uid170: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid170_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid170_Out0_copy171);
   Compressor_6_3_F125_uid69_bh4_uid170_Out0 <= Compressor_6_3_F125_uid69_bh4_uid170_Out0_copy171; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid172_In0 <= "" & bh4_w11_6 & bh4_w11_7 & bh4_w11_0 & bh4_w11_9;
   Compressor_14_3_F125_uid79_bh4_uid172_In1 <= "" & bh4_w12_8;
   bh4_w11_24 <= Compressor_14_3_F125_uid79_bh4_uid172_Out0(0);
   bh4_w12_19 <= Compressor_14_3_F125_uid79_bh4_uid172_Out0(1);
   bh4_w13_14 <= Compressor_14_3_F125_uid79_bh4_uid172_Out0(2);
   Compressor_14_3_F125_uid79_uid172: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid172_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid172_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid172_Out0_copy173);
   Compressor_14_3_F125_uid79_bh4_uid172_Out0 <= Compressor_14_3_F125_uid79_bh4_uid172_Out0_copy173; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid174_In0 <= "" & bh4_w12_10 & bh4_w12_1 & bh4_w12_2 & bh4_w12_3 & bh4_w12_4 & bh4_w12_5;
   bh4_w12_20 <= Compressor_6_3_F125_uid69_bh4_uid174_Out0(0);
   bh4_w13_15 <= Compressor_6_3_F125_uid69_bh4_uid174_Out0(1);
   bh4_w14_10 <= Compressor_6_3_F125_uid69_bh4_uid174_Out0(2);
   Compressor_6_3_F125_uid69_uid174: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid174_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid174_Out0_copy175);
   Compressor_6_3_F125_uid69_bh4_uid174_Out0 <= Compressor_6_3_F125_uid69_bh4_uid174_Out0_copy175; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid176_In0 <= "" & bh4_w12_13 & bh4_w12_12 & bh4_w12_11 & bh4_w12_9 & bh4_w12_0 & bh4_w12_7;
   bh4_w12_21 <= Compressor_6_3_F125_uid69_bh4_uid176_Out0(0);
   bh4_w13_16 <= Compressor_6_3_F125_uid69_bh4_uid176_Out0(1);
   bh4_w14_11 <= Compressor_6_3_F125_uid69_bh4_uid176_Out0(2);
   Compressor_6_3_F125_uid69_uid176: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid176_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid176_Out0_copy177);
   Compressor_6_3_F125_uid69_bh4_uid176_Out0 <= Compressor_6_3_F125_uid69_bh4_uid176_Out0_copy177; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid178_In0 <= "" & bh4_w13_8 & bh4_w13_11 & bh4_w13_10 & bh4_w13_9 & bh4_w13_0 & bh4_w13_7;
   bh4_w13_17 <= Compressor_6_3_F125_uid69_bh4_uid178_Out0(0);
   bh4_w14_12 <= Compressor_6_3_F125_uid69_bh4_uid178_Out0(1);
   bh4_w15_8 <= Compressor_6_3_F125_uid69_bh4_uid178_Out0(2);
   Compressor_6_3_F125_uid69_uid178: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid178_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid178_Out0_copy179);
   Compressor_6_3_F125_uid69_bh4_uid178_Out0 <= Compressor_6_3_F125_uid69_bh4_uid178_Out0_copy179; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid180_In0 <= "" & bh4_w13_1 & bh4_w13_2 & bh4_w13_3 & bh4_w13_4 & bh4_w13_5 & bh4_w13_6;
   bh4_w13_18 <= Compressor_6_3_F125_uid69_bh4_uid180_Out0(0);
   bh4_w14_13 <= Compressor_6_3_F125_uid69_bh4_uid180_Out0(1);
   bh4_w15_9 <= Compressor_6_3_F125_uid69_bh4_uid180_Out0(2);
   Compressor_6_3_F125_uid69_uid180: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid180_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid180_Out0_copy181);
   Compressor_6_3_F125_uid69_bh4_uid180_Out0 <= Compressor_6_3_F125_uid69_bh4_uid180_Out0_copy181; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid182_In0 <= "" & bh4_w14_0 & bh4_w14_1 & bh4_w14_2 & bh4_w14_3 & bh4_w14_4 & bh4_w14_5;
   bh4_w14_14 <= Compressor_6_3_F125_uid69_bh4_uid182_Out0(0);
   bh4_w15_10 <= Compressor_6_3_F125_uid69_bh4_uid182_Out0(1);
   bh4_w16_6 <= Compressor_6_3_F125_uid69_bh4_uid182_Out0(2);
   Compressor_6_3_F125_uid69_uid182: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid182_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid182_Out0_copy183);
   Compressor_6_3_F125_uid69_bh4_uid182_Out0 <= Compressor_6_3_F125_uid69_bh4_uid182_Out0_copy183; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid184_In0 <= "" & bh4_w14_6 & bh4_w14_7 & bh4_w14_8 & bh4_w14_9;
   Compressor_14_3_F125_uid79_bh4_uid184_In1 <= "" & bh4_w15_0;
   bh4_w14_15 <= Compressor_14_3_F125_uid79_bh4_uid184_Out0(0);
   bh4_w15_11 <= Compressor_14_3_F125_uid79_bh4_uid184_Out0(1);
   bh4_w16_7 <= Compressor_14_3_F125_uid79_bh4_uid184_Out0(2);
   Compressor_14_3_F125_uid79_uid184: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid184_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid184_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid184_Out0_copy185);
   Compressor_14_3_F125_uid79_bh4_uid184_Out0 <= Compressor_14_3_F125_uid79_bh4_uid184_Out0_copy185; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid186_In0 <= "" & bh4_w15_1 & bh4_w15_2 & bh4_w15_3 & bh4_w15_4 & bh4_w15_5 & bh4_w15_6;
   bh4_w15_12 <= Compressor_6_3_F125_uid69_bh4_uid186_Out0(0);
   bh4_w16_8 <= Compressor_6_3_F125_uid69_bh4_uid186_Out0(1);
   bh4_w17_5 <= Compressor_6_3_F125_uid69_bh4_uid186_Out0(2);
   Compressor_6_3_F125_uid69_uid186: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid186_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid186_Out0_copy187);
   Compressor_6_3_F125_uid69_bh4_uid186_Out0 <= Compressor_6_3_F125_uid69_bh4_uid186_Out0_copy187; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid188_In0 <= "" & bh4_w16_0 & bh4_w16_1 & bh4_w16_2 & bh4_w16_3 & bh4_w16_4 & bh4_w16_5;
   bh4_w16_9 <= Compressor_6_3_F125_uid69_bh4_uid188_Out0(0);
   bh4_w17_6 <= Compressor_6_3_F125_uid69_bh4_uid188_Out0(1);
   bh4_w18_3 <= Compressor_6_3_F125_uid69_bh4_uid188_Out0(2);
   Compressor_6_3_F125_uid69_uid188: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid188_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid188_Out0_copy189);
   Compressor_6_3_F125_uid69_bh4_uid188_Out0 <= Compressor_6_3_F125_uid69_bh4_uid188_Out0_copy189; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid190_In0 <= "" & bh4_w17_0 & bh4_w17_1 & bh4_w17_2 & bh4_w17_3;
   Compressor_14_3_F125_uid79_bh4_uid190_In1 <= "" & "0";
   bh4_w17_7 <= Compressor_14_3_F125_uid79_bh4_uid190_Out0(0);
   bh4_w18_4 <= Compressor_14_3_F125_uid79_bh4_uid190_Out0(1);
   bh4_w19_2 <= Compressor_14_3_F125_uid79_bh4_uid190_Out0(2);
   Compressor_14_3_F125_uid79_uid190: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid190_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid190_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid190_Out0_copy191);
   Compressor_14_3_F125_uid79_bh4_uid190_Out0 <= Compressor_14_3_F125_uid79_bh4_uid190_Out0_copy191; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid194_In0 <= "" & bh4_w18_0 & bh4_w18_1 & bh4_w18_2;
   Compressor_23_3_F125_uid193_bh4_uid194_In1 <= "" & bh4_w19_0 & bh4_w19_1;
   bh4_w18_5 <= Compressor_23_3_F125_uid193_bh4_uid194_Out0(0);
   bh4_w19_3 <= Compressor_23_3_F125_uid193_bh4_uid194_Out0(1);
   bh4_w20_2 <= Compressor_23_3_F125_uid193_bh4_uid194_Out0(2);
   Compressor_23_3_F125_uid193_uid194: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid194_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid194_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid194_Out0_copy195);
   Compressor_23_3_F125_uid193_bh4_uid194_Out0 <= Compressor_23_3_F125_uid193_bh4_uid194_Out0_copy195; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid196_In0 <= "" & bh4_w20_0 & bh4_w20_1 & "0";
   Compressor_23_3_F125_uid193_bh4_uid196_In1 <= "" & bh4_w21_0 & bh4_w21_1;
   bh4_w20_3 <= Compressor_23_3_F125_uid193_bh4_uid196_Out0(0);
   bh4_w21_2 <= Compressor_23_3_F125_uid193_bh4_uid196_Out0(1);
   bh4_w22_2 <= Compressor_23_3_F125_uid193_bh4_uid196_Out0(2);
   Compressor_23_3_F125_uid193_uid196: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid196_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid196_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid196_Out0_copy197);
   Compressor_23_3_F125_uid193_bh4_uid196_Out0 <= Compressor_23_3_F125_uid193_bh4_uid196_Out0_copy197; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid198_In0 <= "" & bh4_w22_0 & bh4_w22_1 & "0";
   Compressor_23_3_F125_uid193_bh4_uid198_In1 <= "" & bh4_w23_0 & bh4_w23_1;
   bh4_w22_3 <= Compressor_23_3_F125_uid193_bh4_uid198_Out0(0);
   bh4_w23_2 <= Compressor_23_3_F125_uid193_bh4_uid198_Out0(1);
   bh4_w24_2 <= Compressor_23_3_F125_uid193_bh4_uid198_Out0(2);
   Compressor_23_3_F125_uid193_uid198: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid198_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid198_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid198_Out0_copy199);
   Compressor_23_3_F125_uid193_bh4_uid198_Out0 <= Compressor_23_3_F125_uid193_bh4_uid198_Out0_copy199; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid200_In0 <= "" & bh4_w24_0 & bh4_w24_1 & "0";
   Compressor_23_3_F125_uid193_bh4_uid200_In1 <= "" & bh4_w25_0 & bh4_w25_1;
   bh4_w24_3 <= Compressor_23_3_F125_uid193_bh4_uid200_Out0(0);
   bh4_w25_2 <= Compressor_23_3_F125_uid193_bh4_uid200_Out0(1);
   bh4_w26_2 <= Compressor_23_3_F125_uid193_bh4_uid200_Out0(2);
   Compressor_23_3_F125_uid193_uid200: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid200_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid200_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid200_Out0_copy201);
   Compressor_23_3_F125_uid193_bh4_uid200_Out0 <= Compressor_23_3_F125_uid193_bh4_uid200_Out0_copy201; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid202_In0 <= "" & bh4_w26_0 & bh4_w26_1 & "0";
   Compressor_23_3_F125_uid193_bh4_uid202_In1 <= "" & bh4_w27_0 & bh4_w27_1;
   bh4_w26_3 <= Compressor_23_3_F125_uid193_bh4_uid202_Out0(0);
   bh4_w27_2 <= Compressor_23_3_F125_uid193_bh4_uid202_Out0(1);
   bh4_w28_2 <= Compressor_23_3_F125_uid193_bh4_uid202_Out0(2);
   Compressor_23_3_F125_uid193_uid202: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid202_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid202_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid202_Out0_copy203);
   Compressor_23_3_F125_uid193_bh4_uid202_Out0 <= Compressor_23_3_F125_uid193_bh4_uid202_Out0_copy203; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid204_In0 <= "" & bh4_w28_0 & bh4_w28_1 & "0";
   Compressor_23_3_F125_uid193_bh4_uid204_In1 <= "" & bh4_w29_0 & bh4_w29_1;
   bh4_w28_3 <= Compressor_23_3_F125_uid193_bh4_uid204_Out0(0);
   bh4_w29_2 <= Compressor_23_3_F125_uid193_bh4_uid204_Out0(1);
   bh4_w30_2 <= Compressor_23_3_F125_uid193_bh4_uid204_Out0(2);
   Compressor_23_3_F125_uid193_uid204: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid204_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid204_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid204_Out0_copy205);
   Compressor_23_3_F125_uid193_bh4_uid204_Out0 <= Compressor_23_3_F125_uid193_bh4_uid204_Out0_copy205; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid206_In0 <= "" & bh4_w30_0 & bh4_w30_1 & "0";
   Compressor_23_3_F125_uid193_bh4_uid206_In1 <= "" & bh4_w31_0 & bh4_w31_1;
   bh4_w30_3 <= Compressor_23_3_F125_uid193_bh4_uid206_Out0(0);
   bh4_w31_2 <= Compressor_23_3_F125_uid193_bh4_uid206_Out0(1);
   bh4_w32_2 <= Compressor_23_3_F125_uid193_bh4_uid206_Out0(2);
   Compressor_23_3_F125_uid193_uid206: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid206_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid206_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid206_Out0_copy207);
   Compressor_23_3_F125_uid193_bh4_uid206_Out0 <= Compressor_23_3_F125_uid193_bh4_uid206_Out0_copy207; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid208_In0 <= "" & bh4_w32_0 & bh4_w32_1 & "0";
   Compressor_23_3_F125_uid193_bh4_uid208_In1 <= "" & bh4_w33_0 & bh4_w33_1;
   bh4_w32_3 <= Compressor_23_3_F125_uid193_bh4_uid208_Out0(0);
   bh4_w33_2 <= Compressor_23_3_F125_uid193_bh4_uid208_Out0(1);
   bh4_w34_2 <= Compressor_23_3_F125_uid193_bh4_uid208_Out0(2);
   Compressor_23_3_F125_uid193_uid208: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid208_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid208_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid208_Out0_copy209);
   Compressor_23_3_F125_uid193_bh4_uid208_Out0 <= Compressor_23_3_F125_uid193_bh4_uid208_Out0_copy209; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid210_In0 <= "" & bh4_w34_0 & bh4_w34_1 & "0";
   Compressor_23_3_F125_uid193_bh4_uid210_In1 <= "" & bh4_w35_0 & bh4_w35_1;
   bh4_w34_3 <= Compressor_23_3_F125_uid193_bh4_uid210_Out0(0);
   bh4_w35_2 <= Compressor_23_3_F125_uid193_bh4_uid210_Out0(1);
   bh4_w36_1 <= Compressor_23_3_F125_uid193_bh4_uid210_Out0(2);
   Compressor_23_3_F125_uid193_uid210: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid210_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid210_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid210_Out0_copy211);
   Compressor_23_3_F125_uid193_bh4_uid210_Out0 <= Compressor_23_3_F125_uid193_bh4_uid210_Out0_copy211; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid212_In0 <= "" & bh4_w0_33 & bh4_w0_31 & bh4_w0_29 & bh4_w0_30 & bh4_w0_32 & bh4_w0_12;
   bh4_w0_34 <= Compressor_6_3_F125_uid69_bh4_uid212_Out0(0);
   bh4_w1_41 <= Compressor_6_3_F125_uid69_bh4_uid212_Out0(1);
   bh4_w2_46 <= Compressor_6_3_F125_uid69_bh4_uid212_Out0(2);
   Compressor_6_3_F125_uid69_uid212: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid212_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid212_Out0_copy213);
   Compressor_6_3_F125_uid69_bh4_uid212_Out0 <= Compressor_6_3_F125_uid69_bh4_uid212_Out0_copy213; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid214_In0 <= "" & bh4_w1_36 & bh4_w1_34 & bh4_w1_33 & bh4_w1_31 & bh4_w1_32 & bh4_w1_39;
   bh4_w1_42 <= Compressor_6_3_F125_uid69_bh4_uid214_Out0(0);
   bh4_w2_47 <= Compressor_6_3_F125_uid69_bh4_uid214_Out0(1);
   bh4_w3_46 <= Compressor_6_3_F125_uid69_bh4_uid214_Out0(2);
   Compressor_6_3_F125_uid69_uid214: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid214_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid214_Out0_copy215);
   Compressor_6_3_F125_uid69_bh4_uid214_Out0 <= Compressor_6_3_F125_uid69_bh4_uid214_Out0_copy215; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid216_In0 <= "" & bh4_w1_37 & bh4_w1_35 & bh4_w1_40 & bh4_w1_38;
   Compressor_14_3_F125_uid79_bh4_uid216_In1 <= "" & bh4_w2_37;
   bh4_w1_43 <= Compressor_14_3_F125_uid79_bh4_uid216_Out0(0);
   bh4_w2_48 <= Compressor_14_3_F125_uid79_bh4_uid216_Out0(1);
   bh4_w3_47 <= Compressor_14_3_F125_uid79_bh4_uid216_Out0(2);
   Compressor_14_3_F125_uid79_uid216: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid216_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid216_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid216_Out0_copy217);
   Compressor_14_3_F125_uid79_bh4_uid216_Out0 <= Compressor_14_3_F125_uid79_bh4_uid216_Out0_copy217; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid218_In0 <= "" & bh4_w2_1 & bh4_w2_39 & bh4_w2_32 & bh4_w2_31 & bh4_w2_33 & bh4_w2_34;
   bh4_w2_49 <= Compressor_6_3_F125_uid69_bh4_uid218_Out0(0);
   bh4_w3_48 <= Compressor_6_3_F125_uid69_bh4_uid218_Out0(1);
   bh4_w4_46 <= Compressor_6_3_F125_uid69_bh4_uid218_Out0(2);
   Compressor_6_3_F125_uid69_uid218: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid218_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid218_Out0_copy219);
   Compressor_6_3_F125_uid69_bh4_uid218_Out0 <= Compressor_6_3_F125_uid69_bh4_uid218_Out0_copy219; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid220_In0 <= "" & bh4_w2_44 & bh4_w2_42 & bh4_w2_40 & bh4_w2_45 & bh4_w2_43 & bh4_w2_41;
   bh4_w2_50 <= Compressor_6_3_F125_uid69_bh4_uid220_Out0(0);
   bh4_w3_49 <= Compressor_6_3_F125_uid69_bh4_uid220_Out0(1);
   bh4_w4_47 <= Compressor_6_3_F125_uid69_bh4_uid220_Out0(2);
   Compressor_6_3_F125_uid69_uid220: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid220_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid220_Out0_copy221);
   Compressor_6_3_F125_uid69_bh4_uid220_Out0 <= Compressor_6_3_F125_uid69_bh4_uid220_Out0_copy221; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid224_In0 <= "" & bh4_w2_36 & bh4_w2_38 & bh4_w2_35;
   bh4_w2_51 <= Compressor_3_2_F125_uid223_bh4_uid224_Out0(0);
   bh4_w3_50 <= Compressor_3_2_F125_uid223_bh4_uid224_Out0(1);
   Compressor_3_2_F125_uid223_uid224: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid224_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid224_Out0_copy225);
   Compressor_3_2_F125_uid223_bh4_uid224_Out0 <= Compressor_3_2_F125_uid223_bh4_uid224_Out0_copy225; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid226_In0 <= "" & bh4_w3_36 & bh4_w3_40 & bh4_w3_42 & bh4_w3_44 & bh4_w3_30 & bh4_w3_32;
   bh4_w3_51 <= Compressor_6_3_F125_uid69_bh4_uid226_Out0(0);
   bh4_w4_48 <= Compressor_6_3_F125_uid69_bh4_uid226_Out0(1);
   bh4_w5_43 <= Compressor_6_3_F125_uid69_bh4_uid226_Out0(2);
   Compressor_6_3_F125_uid69_uid226: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid226_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid226_Out0_copy227);
   Compressor_6_3_F125_uid69_bh4_uid226_Out0 <= Compressor_6_3_F125_uid69_bh4_uid226_Out0_copy227; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid228_In0 <= "" & bh4_w3_34 & bh4_w3_45 & bh4_w3_43 & bh4_w3_41 & bh4_w3_39 & bh4_w3_37;
   bh4_w3_52 <= Compressor_6_3_F125_uid69_bh4_uid228_Out0(0);
   bh4_w4_49 <= Compressor_6_3_F125_uid69_bh4_uid228_Out0(1);
   bh4_w5_44 <= Compressor_6_3_F125_uid69_bh4_uid228_Out0(2);
   Compressor_6_3_F125_uid69_uid228: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid228_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid228_Out0_copy229);
   Compressor_6_3_F125_uid69_bh4_uid228_Out0 <= Compressor_6_3_F125_uid69_bh4_uid228_Out0_copy229; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid230_In0 <= "" & bh4_w3_31 & bh4_w3_33 & bh4_w3_38 & bh4_w3_35;
   Compressor_14_3_F125_uid79_bh4_uid230_In1 <= "" & bh4_w4_37;
   bh4_w3_53 <= Compressor_14_3_F125_uid79_bh4_uid230_Out0(0);
   bh4_w4_50 <= Compressor_14_3_F125_uid79_bh4_uid230_Out0(1);
   bh4_w5_45 <= Compressor_14_3_F125_uid79_bh4_uid230_Out0(2);
   Compressor_14_3_F125_uid79_uid230: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid230_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid230_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid230_Out0_copy231);
   Compressor_14_3_F125_uid79_bh4_uid230_Out0 <= Compressor_14_3_F125_uid79_bh4_uid230_Out0_copy231; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid232_In0 <= "" & bh4_w4_35 & bh4_w4_44 & bh4_w4_42 & bh4_w4_40 & bh4_w4_45 & bh4_w4_43;
   bh4_w4_51 <= Compressor_6_3_F125_uid69_bh4_uid232_Out0(0);
   bh4_w5_46 <= Compressor_6_3_F125_uid69_bh4_uid232_Out0(1);
   bh4_w6_40 <= Compressor_6_3_F125_uid69_bh4_uid232_Out0(2);
   Compressor_6_3_F125_uid69_uid232: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid232_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid232_Out0_copy233);
   Compressor_6_3_F125_uid69_bh4_uid232_Out0 <= Compressor_6_3_F125_uid69_bh4_uid232_Out0_copy233; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid234_In0 <= "" & bh4_w4_39 & bh4_w4_32 & bh4_w4_31 & bh4_w4_33 & bh4_w4_34 & bh4_w4_36;
   bh4_w4_52 <= Compressor_6_3_F125_uid69_bh4_uid234_Out0(0);
   bh4_w5_47 <= Compressor_6_3_F125_uid69_bh4_uid234_Out0(1);
   bh4_w6_41 <= Compressor_6_3_F125_uid69_bh4_uid234_Out0(2);
   Compressor_6_3_F125_uid69_uid234: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid234_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid234_Out0_copy235);
   Compressor_6_3_F125_uid69_bh4_uid234_Out0 <= Compressor_6_3_F125_uid69_bh4_uid234_Out0_copy235; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid236_In0 <= "" & bh4_w4_41 & bh4_w4_1 & bh4_w4_38;
   Compressor_23_3_F125_uid193_bh4_uid236_In1 <= "" & bh4_w5_38 & bh4_w5_41;
   bh4_w4_53 <= Compressor_23_3_F125_uid193_bh4_uid236_Out0(0);
   bh4_w5_48 <= Compressor_23_3_F125_uid193_bh4_uid236_Out0(1);
   bh4_w6_42 <= Compressor_23_3_F125_uid193_bh4_uid236_Out0(2);
   Compressor_23_3_F125_uid193_uid236: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid236_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid236_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid236_Out0_copy237);
   Compressor_23_3_F125_uid193_bh4_uid236_Out0 <= Compressor_23_3_F125_uid193_bh4_uid236_Out0_copy237; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid238_In0 <= "" & bh4_w5_40 & bh4_w5_31 & bh4_w5_29 & bh4_w5_28 & bh4_w5_30 & bh4_w5_32;
   bh4_w5_49 <= Compressor_6_3_F125_uid69_bh4_uid238_Out0(0);
   bh4_w6_43 <= Compressor_6_3_F125_uid69_bh4_uid238_Out0(1);
   bh4_w7_37 <= Compressor_6_3_F125_uid69_bh4_uid238_Out0(2);
   Compressor_6_3_F125_uid69_uid238: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid238_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid238_Out0_copy239);
   Compressor_6_3_F125_uid69_bh4_uid238_Out0 <= Compressor_6_3_F125_uid69_bh4_uid238_Out0_copy239; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid240_In0 <= "" & bh4_w5_39 & bh4_w5_37 & bh4_w5_35 & bh4_w5_33 & bh4_w5_42 & bh4_w5_36;
   bh4_w5_50 <= Compressor_6_3_F125_uid69_bh4_uid240_Out0(0);
   bh4_w6_44 <= Compressor_6_3_F125_uid69_bh4_uid240_Out0(1);
   bh4_w7_38 <= Compressor_6_3_F125_uid69_bh4_uid240_Out0(2);
   Compressor_6_3_F125_uid69_uid240: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid240_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid240_Out0_copy241);
   Compressor_6_3_F125_uid69_bh4_uid240_Out0 <= Compressor_6_3_F125_uid69_bh4_uid240_Out0_copy241; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid242_In0 <= "" & bh4_w6_26 & bh4_w6_39 & bh4_w6_37 & bh4_w6_35 & bh4_w6_33 & bh4_w6_32;
   bh4_w6_45 <= Compressor_6_3_F125_uid69_bh4_uid242_Out0(0);
   bh4_w7_39 <= Compressor_6_3_F125_uid69_bh4_uid242_Out0(1);
   bh4_w8_34 <= Compressor_6_3_F125_uid69_bh4_uid242_Out0(2);
   Compressor_6_3_F125_uid69_uid242: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid242_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid242_Out0_copy243);
   Compressor_6_3_F125_uid69_bh4_uid242_Out0 <= Compressor_6_3_F125_uid69_bh4_uid242_Out0_copy243; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid244_In0 <= "" & bh4_w6_28 & bh4_w6_22 & bh4_w6_31 & bh4_w6_29 & bh4_w6_27 & bh4_w6_34;
   bh4_w6_46 <= Compressor_6_3_F125_uid69_bh4_uid244_Out0(0);
   bh4_w7_40 <= Compressor_6_3_F125_uid69_bh4_uid244_Out0(1);
   bh4_w8_35 <= Compressor_6_3_F125_uid69_bh4_uid244_Out0(2);
   Compressor_6_3_F125_uid69_uid244: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid244_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid244_Out0_copy245);
   Compressor_6_3_F125_uid69_bh4_uid244_Out0 <= Compressor_6_3_F125_uid69_bh4_uid244_Out0_copy245; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid246_In0 <= "" & bh4_w6_30 & bh4_w6_38 & bh4_w6_36;
   bh4_w6_47 <= Compressor_3_2_F125_uid223_bh4_uid246_Out0(0);
   bh4_w7_41 <= Compressor_3_2_F125_uid223_bh4_uid246_Out0(1);
   Compressor_3_2_F125_uid223_uid246: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid246_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid246_Out0_copy247);
   Compressor_3_2_F125_uid223_bh4_uid246_Out0 <= Compressor_3_2_F125_uid223_bh4_uid246_Out0_copy247; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid248_In0 <= "" & bh4_w7_35 & bh4_w7_36 & bh4_w7_34 & bh4_w7_31 & bh4_w7_32 & bh4_w7_33;
   bh4_w7_42 <= Compressor_6_3_F125_uid69_bh4_uid248_Out0(0);
   bh4_w8_36 <= Compressor_6_3_F125_uid69_bh4_uid248_Out0(1);
   bh4_w9_31 <= Compressor_6_3_F125_uid69_bh4_uid248_Out0(2);
   Compressor_6_3_F125_uid69_uid248: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid248_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid248_Out0_copy249);
   Compressor_6_3_F125_uid69_bh4_uid248_Out0 <= Compressor_6_3_F125_uid69_bh4_uid248_Out0_copy249; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid250_In0 <= "" & bh4_w7_30 & bh4_w7_29 & bh4_w7_27 & bh4_w7_25 & bh4_w7_24 & bh4_w7_26;
   bh4_w7_43 <= Compressor_6_3_F125_uid69_bh4_uid250_Out0(0);
   bh4_w8_37 <= Compressor_6_3_F125_uid69_bh4_uid250_Out0(1);
   bh4_w9_32 <= Compressor_6_3_F125_uid69_bh4_uid250_Out0(2);
   Compressor_6_3_F125_uid69_uid250: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid250_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid250_Out0_copy251);
   Compressor_6_3_F125_uid69_bh4_uid250_Out0 <= Compressor_6_3_F125_uid69_bh4_uid250_Out0_copy251; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid252_In0 <= "" & bh4_w8_33 & bh4_w8_26 & bh4_w8_32 & bh4_w8_30 & bh4_w8_28 & bh4_w8_24;
   bh4_w8_38 <= Compressor_6_3_F125_uid69_bh4_uid252_Out0(0);
   bh4_w9_33 <= Compressor_6_3_F125_uid69_bh4_uid252_Out0(1);
   bh4_w10_28 <= Compressor_6_3_F125_uid69_bh4_uid252_Out0(2);
   Compressor_6_3_F125_uid69_uid252: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid252_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid252_Out0_copy253);
   Compressor_6_3_F125_uid69_bh4_uid252_Out0 <= Compressor_6_3_F125_uid69_bh4_uid252_Out0_copy253; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid254_In0 <= "" & bh4_w8_31 & bh4_w8_29 & bh4_w8_27 & bh4_w8_25 & bh4_w8_23 & bh4_w8_22;
   bh4_w8_39 <= Compressor_6_3_F125_uid69_bh4_uid254_Out0(0);
   bh4_w9_34 <= Compressor_6_3_F125_uid69_bh4_uid254_Out0(1);
   bh4_w10_29 <= Compressor_6_3_F125_uid69_bh4_uid254_Out0(2);
   Compressor_6_3_F125_uid69_uid254: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid254_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid254_Out0_copy255);
   Compressor_6_3_F125_uid69_bh4_uid254_Out0 <= Compressor_6_3_F125_uid69_bh4_uid254_Out0_copy255; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid256_In0 <= "" & bh4_w9_29 & bh4_w9_27 & bh4_w9_25 & bh4_w9_23 & bh4_w9_21 & bh4_w9_20;
   bh4_w9_35 <= Compressor_6_3_F125_uid69_bh4_uid256_Out0(0);
   bh4_w10_30 <= Compressor_6_3_F125_uid69_bh4_uid256_Out0(1);
   bh4_w11_25 <= Compressor_6_3_F125_uid69_bh4_uid256_Out0(2);
   Compressor_6_3_F125_uid69_uid256: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid256_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid256_Out0_copy257);
   Compressor_6_3_F125_uid69_bh4_uid256_Out0 <= Compressor_6_3_F125_uid69_bh4_uid256_Out0_copy257; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid258_In0 <= "" & bh4_w9_8 & bh4_w9_30 & bh4_w9_28 & bh4_w9_26 & bh4_w9_24 & bh4_w9_22;
   bh4_w9_36 <= Compressor_6_3_F125_uid69_bh4_uid258_Out0(0);
   bh4_w10_31 <= Compressor_6_3_F125_uid69_bh4_uid258_Out0(1);
   bh4_w11_26 <= Compressor_6_3_F125_uid69_bh4_uid258_Out0(2);
   Compressor_6_3_F125_uid69_uid258: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid258_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid258_Out0_copy259);
   Compressor_6_3_F125_uid69_bh4_uid258_Out0 <= Compressor_6_3_F125_uid69_bh4_uid258_Out0_copy259; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid260_In0 <= "" & bh4_w10_27 & bh4_w10_25 & bh4_w10_23 & bh4_w10_21 & bh4_w10_19 & bh4_w10_18;
   bh4_w10_32 <= Compressor_6_3_F125_uid69_bh4_uid260_Out0(0);
   bh4_w11_27 <= Compressor_6_3_F125_uid69_bh4_uid260_Out0(1);
   bh4_w12_22 <= Compressor_6_3_F125_uid69_bh4_uid260_Out0(2);
   Compressor_6_3_F125_uid69_uid260: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid260_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid260_Out0_copy261);
   Compressor_6_3_F125_uid69_bh4_uid260_Out0 <= Compressor_6_3_F125_uid69_bh4_uid260_Out0_copy261; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid262_In0 <= "" & bh4_w10_20 & bh4_w10_22 & bh4_w10_24 & bh4_w10_26;
   Compressor_14_3_F125_uid79_bh4_uid262_In1 <= "" & "0";
   bh4_w10_33 <= Compressor_14_3_F125_uid79_bh4_uid262_Out0(0);
   bh4_w11_28 <= Compressor_14_3_F125_uid79_bh4_uid262_Out0(1);
   bh4_w12_23 <= Compressor_14_3_F125_uid79_bh4_uid262_Out0(2);
   Compressor_14_3_F125_uid79_uid262: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid262_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid262_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid262_Out0_copy263);
   Compressor_14_3_F125_uid79_bh4_uid262_Out0 <= Compressor_14_3_F125_uid79_bh4_uid262_Out0_copy263; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid264_In0 <= "" & bh4_w11_23 & bh4_w11_21 & bh4_w11_19 & bh4_w11_17 & bh4_w11_16 & bh4_w11_18;
   bh4_w11_29 <= Compressor_6_3_F125_uid69_bh4_uid264_Out0(0);
   bh4_w12_24 <= Compressor_6_3_F125_uid69_bh4_uid264_Out0(1);
   bh4_w13_19 <= Compressor_6_3_F125_uid69_bh4_uid264_Out0(2);
   Compressor_6_3_F125_uid69_uid264: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid264_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid264_Out0_copy265);
   Compressor_6_3_F125_uid69_bh4_uid264_Out0 <= Compressor_6_3_F125_uid69_bh4_uid264_Out0_copy265; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid266_In0 <= "" & bh4_w11_20 & bh4_w11_22 & bh4_w11_24;
   bh4_w11_30 <= Compressor_3_2_F125_uid223_bh4_uid266_Out0(0);
   bh4_w12_25 <= Compressor_3_2_F125_uid223_bh4_uid266_Out0(1);
   Compressor_3_2_F125_uid223_uid266: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid266_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid266_Out0_copy267);
   Compressor_3_2_F125_uid223_bh4_uid266_Out0 <= Compressor_3_2_F125_uid223_bh4_uid266_Out0_copy267; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid268_In0 <= "" & bh4_w12_6 & bh4_w12_20 & bh4_w12_18 & bh4_w12_16 & bh4_w12_15 & bh4_w12_14;
   bh4_w12_26 <= Compressor_6_3_F125_uid69_bh4_uid268_Out0(0);
   bh4_w13_20 <= Compressor_6_3_F125_uid69_bh4_uid268_Out0(1);
   bh4_w14_16 <= Compressor_6_3_F125_uid69_bh4_uid268_Out0(2);
   Compressor_6_3_F125_uid69_uid268: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid268_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid268_Out0_copy269);
   Compressor_6_3_F125_uid69_bh4_uid268_Out0 <= Compressor_6_3_F125_uid69_bh4_uid268_Out0_copy269; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid270_In0 <= "" & bh4_w12_17 & bh4_w12_19 & bh4_w12_21;
   bh4_w12_27 <= Compressor_3_2_F125_uid223_bh4_uid270_Out0(0);
   bh4_w13_21 <= Compressor_3_2_F125_uid223_bh4_uid270_Out0(1);
   Compressor_3_2_F125_uid223_uid270: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid270_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid270_Out0_copy271);
   Compressor_3_2_F125_uid223_bh4_uid270_Out0 <= Compressor_3_2_F125_uid223_bh4_uid270_Out0_copy271; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid272_In0 <= "" & bh4_w13_17 & bh4_w13_12 & bh4_w13_13 & bh4_w13_14 & bh4_w13_15 & bh4_w13_16;
   bh4_w13_22 <= Compressor_6_3_F125_uid69_bh4_uid272_Out0(0);
   bh4_w14_17 <= Compressor_6_3_F125_uid69_bh4_uid272_Out0(1);
   bh4_w15_13 <= Compressor_6_3_F125_uid69_bh4_uid272_Out0(2);
   Compressor_6_3_F125_uid69_uid272: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid272_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid272_Out0_copy273);
   Compressor_6_3_F125_uid69_bh4_uid272_Out0 <= Compressor_6_3_F125_uid69_bh4_uid272_Out0_copy273; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid274_In0 <= "" & bh4_w14_15 & bh4_w14_14 & bh4_w14_13 & bh4_w14_12 & bh4_w14_11 & bh4_w14_10;
   bh4_w14_18 <= Compressor_6_3_F125_uid69_bh4_uid274_Out0(0);
   bh4_w15_14 <= Compressor_6_3_F125_uid69_bh4_uid274_Out0(1);
   bh4_w16_10 <= Compressor_6_3_F125_uid69_bh4_uid274_Out0(2);
   Compressor_6_3_F125_uid69_uid274: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid274_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid274_Out0_copy275);
   Compressor_6_3_F125_uid69_bh4_uid274_Out0 <= Compressor_6_3_F125_uid69_bh4_uid274_Out0_copy275; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid276_In0 <= "" & bh4_w15_7 & bh4_w15_12 & bh4_w15_11 & bh4_w15_10 & bh4_w15_9 & bh4_w15_8;
   bh4_w15_15 <= Compressor_6_3_F125_uid69_bh4_uid276_Out0(0);
   bh4_w16_11 <= Compressor_6_3_F125_uid69_bh4_uid276_Out0(1);
   bh4_w17_8 <= Compressor_6_3_F125_uid69_bh4_uid276_Out0(2);
   Compressor_6_3_F125_uid69_uid276: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid276_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid276_Out0_copy277);
   Compressor_6_3_F125_uid69_bh4_uid276_Out0 <= Compressor_6_3_F125_uid69_bh4_uid276_Out0_copy277; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid278_In0 <= "" & bh4_w16_9 & bh4_w16_8 & bh4_w16_7 & bh4_w16_6;
   Compressor_14_3_F125_uid79_bh4_uid278_In1 <= "" & bh4_w17_4;
   bh4_w16_12 <= Compressor_14_3_F125_uid79_bh4_uid278_Out0(0);
   bh4_w17_9 <= Compressor_14_3_F125_uid79_bh4_uid278_Out0(1);
   bh4_w18_6 <= Compressor_14_3_F125_uid79_bh4_uid278_Out0(2);
   Compressor_14_3_F125_uid79_uid278: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid278_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid278_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid278_Out0_copy279);
   Compressor_14_3_F125_uid79_bh4_uid278_Out0 <= Compressor_14_3_F125_uid79_bh4_uid278_Out0_copy279; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid280_In0 <= "" & bh4_w17_7 & bh4_w17_6 & bh4_w17_5;
   Compressor_23_3_F125_uid193_bh4_uid280_In1 <= "" & bh4_w18_5 & bh4_w18_4;
   bh4_w17_10 <= Compressor_23_3_F125_uid193_bh4_uid280_Out0(0);
   bh4_w18_7 <= Compressor_23_3_F125_uid193_bh4_uid280_Out0(1);
   bh4_w19_4 <= Compressor_23_3_F125_uid193_bh4_uid280_Out0(2);
   Compressor_23_3_F125_uid193_uid280: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid280_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid280_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid280_Out0_copy281);
   Compressor_23_3_F125_uid193_bh4_uid280_Out0 <= Compressor_23_3_F125_uid193_bh4_uid280_Out0_copy281; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid282_In0 <= "" & bh4_w19_3 & bh4_w19_2 & "0";
   Compressor_23_3_F125_uid193_bh4_uid282_In1 <= "" & bh4_w20_3 & bh4_w20_2;
   bh4_w19_5 <= Compressor_23_3_F125_uid193_bh4_uid282_Out0(0);
   bh4_w20_4 <= Compressor_23_3_F125_uid193_bh4_uid282_Out0(1);
   bh4_w21_3 <= Compressor_23_3_F125_uid193_bh4_uid282_Out0(2);
   Compressor_23_3_F125_uid193_uid282: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid282_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid282_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid282_Out0_copy283);
   Compressor_23_3_F125_uid193_bh4_uid282_Out0 <= Compressor_23_3_F125_uid193_bh4_uid282_Out0_copy283; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid284_In0 <= "" & bh4_w22_3 & bh4_w22_2 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid284_In1 <= "" & bh4_w23_2;
   bh4_w22_4 <= Compressor_14_3_F125_uid79_bh4_uid284_Out0(0);
   bh4_w23_3 <= Compressor_14_3_F125_uid79_bh4_uid284_Out0(1);
   bh4_w24_4 <= Compressor_14_3_F125_uid79_bh4_uid284_Out0(2);
   Compressor_14_3_F125_uid79_uid284: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid284_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid284_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid284_Out0_copy285);
   Compressor_14_3_F125_uid79_bh4_uid284_Out0 <= Compressor_14_3_F125_uid79_bh4_uid284_Out0_copy285; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid286_In0 <= "" & bh4_w24_3 & bh4_w24_2 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid286_In1 <= "" & bh4_w25_2;
   bh4_w24_5 <= Compressor_14_3_F125_uid79_bh4_uid286_Out0(0);
   bh4_w25_3 <= Compressor_14_3_F125_uid79_bh4_uid286_Out0(1);
   bh4_w26_4 <= Compressor_14_3_F125_uid79_bh4_uid286_Out0(2);
   Compressor_14_3_F125_uid79_uid286: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid286_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid286_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid286_Out0_copy287);
   Compressor_14_3_F125_uid79_bh4_uid286_Out0 <= Compressor_14_3_F125_uid79_bh4_uid286_Out0_copy287; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid288_In0 <= "" & bh4_w26_3 & bh4_w26_2 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid288_In1 <= "" & bh4_w27_2;
   bh4_w26_5 <= Compressor_14_3_F125_uid79_bh4_uid288_Out0(0);
   bh4_w27_3 <= Compressor_14_3_F125_uid79_bh4_uid288_Out0(1);
   bh4_w28_4 <= Compressor_14_3_F125_uid79_bh4_uid288_Out0(2);
   Compressor_14_3_F125_uid79_uid288: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid288_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid288_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid288_Out0_copy289);
   Compressor_14_3_F125_uid79_bh4_uid288_Out0 <= Compressor_14_3_F125_uid79_bh4_uid288_Out0_copy289; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid290_In0 <= "" & bh4_w28_3 & bh4_w28_2 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid290_In1 <= "" & bh4_w29_2;
   bh4_w28_5 <= Compressor_14_3_F125_uid79_bh4_uid290_Out0(0);
   bh4_w29_3 <= Compressor_14_3_F125_uid79_bh4_uid290_Out0(1);
   bh4_w30_4 <= Compressor_14_3_F125_uid79_bh4_uid290_Out0(2);
   Compressor_14_3_F125_uid79_uid290: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid290_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid290_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid290_Out0_copy291);
   Compressor_14_3_F125_uid79_bh4_uid290_Out0 <= Compressor_14_3_F125_uid79_bh4_uid290_Out0_copy291; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid292_In0 <= "" & bh4_w30_3 & bh4_w30_2 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid292_In1 <= "" & bh4_w31_2;
   bh4_w30_5 <= Compressor_14_3_F125_uid79_bh4_uid292_Out0(0);
   bh4_w31_3 <= Compressor_14_3_F125_uid79_bh4_uid292_Out0(1);
   bh4_w32_4 <= Compressor_14_3_F125_uid79_bh4_uid292_Out0(2);
   Compressor_14_3_F125_uid79_uid292: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid292_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid292_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid292_Out0_copy293);
   Compressor_14_3_F125_uid79_bh4_uid292_Out0 <= Compressor_14_3_F125_uid79_bh4_uid292_Out0_copy293; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid294_In0 <= "" & bh4_w32_3 & bh4_w32_2 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid294_In1 <= "" & bh4_w33_2;
   bh4_w32_5 <= Compressor_14_3_F125_uid79_bh4_uid294_Out0(0);
   bh4_w33_3 <= Compressor_14_3_F125_uid79_bh4_uid294_Out0(1);
   bh4_w34_4 <= Compressor_14_3_F125_uid79_bh4_uid294_Out0(2);
   Compressor_14_3_F125_uid79_uid294: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid294_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid294_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid294_Out0_copy295);
   Compressor_14_3_F125_uid79_bh4_uid294_Out0 <= Compressor_14_3_F125_uid79_bh4_uid294_Out0_copy295; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid296_In0 <= "" & bh4_w34_3 & bh4_w34_2 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid296_In1 <= "" & bh4_w35_2;
   bh4_w34_5 <= Compressor_14_3_F125_uid79_bh4_uid296_Out0(0);
   bh4_w35_3 <= Compressor_14_3_F125_uid79_bh4_uid296_Out0(1);
   bh4_w36_2 <= Compressor_14_3_F125_uid79_bh4_uid296_Out0(2);
   Compressor_14_3_F125_uid79_uid296: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid296_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid296_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid296_Out0_copy297);
   Compressor_14_3_F125_uid79_bh4_uid296_Out0 <= Compressor_14_3_F125_uid79_bh4_uid296_Out0_copy297; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid298_In0 <= "" & bh4_w36_0 & bh4_w36_1 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid298_In1 <= "" & bh4_w37_0;
   bh4_w36_3 <= Compressor_14_3_F125_uid79_bh4_uid298_Out0(0);
   bh4_w37_1 <= Compressor_14_3_F125_uid79_bh4_uid298_Out0(1);
   bh4_w38_1 <= Compressor_14_3_F125_uid79_bh4_uid298_Out0(2);
   Compressor_14_3_F125_uid79_uid298: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid298_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid298_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid298_Out0_copy299);
   Compressor_14_3_F125_uid79_bh4_uid298_Out0 <= Compressor_14_3_F125_uid79_bh4_uid298_Out0_copy299; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid300_In0 <= "" & bh4_w1_43 & bh4_w1_42 & bh4_w1_41;
   bh4_w1_44 <= Compressor_3_2_F125_uid223_bh4_uid300_Out0(0);
   bh4_w2_52 <= Compressor_3_2_F125_uid223_bh4_uid300_Out0(1);
   Compressor_3_2_F125_uid223_uid300: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid300_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid300_Out0_copy301);
   Compressor_3_2_F125_uid223_bh4_uid300_Out0 <= Compressor_3_2_F125_uid223_bh4_uid300_Out0_copy301; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid302_In0 <= "" & bh4_w2_51 & bh4_w2_48 & bh4_w2_49 & bh4_w2_50 & bh4_w2_46 & bh4_w2_47;
   bh4_w2_53 <= Compressor_6_3_F125_uid69_bh4_uid302_Out0(0);
   bh4_w3_54 <= Compressor_6_3_F125_uid69_bh4_uid302_Out0(1);
   bh4_w4_54 <= Compressor_6_3_F125_uid69_bh4_uid302_Out0(2);
   Compressor_6_3_F125_uid69_uid302: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid302_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid302_Out0_copy303);
   Compressor_6_3_F125_uid69_bh4_uid302_Out0 <= Compressor_6_3_F125_uid69_bh4_uid302_Out0_copy303; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid304_In0 <= "" & bh4_w3_51 & bh4_w3_49 & bh4_w3_47 & bh4_w3_52 & bh4_w3_53 & "0";
   bh4_w3_55 <= Compressor_6_3_F125_uid69_bh4_uid304_Out0(0);
   bh4_w4_55 <= Compressor_6_3_F125_uid69_bh4_uid304_Out0(1);
   bh4_w5_51 <= Compressor_6_3_F125_uid69_bh4_uid304_Out0(2);
   Compressor_6_3_F125_uid69_uid304: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid304_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid304_Out0_copy305);
   Compressor_6_3_F125_uid69_bh4_uid304_Out0 <= Compressor_6_3_F125_uid69_bh4_uid304_Out0_copy305; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid306_In0 <= "" & bh4_w3_46 & bh4_w3_48 & bh4_w3_50;
   Compressor_23_3_F125_uid193_bh4_uid306_In1 <= "" & bh4_w4_53 & bh4_w4_50;
   bh4_w3_56 <= Compressor_23_3_F125_uid193_bh4_uid306_Out0(0);
   bh4_w4_56 <= Compressor_23_3_F125_uid193_bh4_uid306_Out0(1);
   bh4_w5_52 <= Compressor_23_3_F125_uid193_bh4_uid306_Out0(2);
   Compressor_23_3_F125_uid193_uid306: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid306_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid306_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid306_Out0_copy307);
   Compressor_23_3_F125_uid193_bh4_uid306_Out0 <= Compressor_23_3_F125_uid193_bh4_uid306_Out0_copy307; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid308_In0 <= "" & bh4_w4_48 & bh4_w4_46 & bh4_w4_51 & bh4_w4_52 & bh4_w4_47 & bh4_w4_49;
   bh4_w4_57 <= Compressor_6_3_F125_uid69_bh4_uid308_Out0(0);
   bh4_w5_53 <= Compressor_6_3_F125_uid69_bh4_uid308_Out0(1);
   bh4_w6_48 <= Compressor_6_3_F125_uid69_bh4_uid308_Out0(2);
   Compressor_6_3_F125_uid69_uid308: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid308_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid308_Out0_copy309);
   Compressor_6_3_F125_uid69_bh4_uid308_Out0 <= Compressor_6_3_F125_uid69_bh4_uid308_Out0_copy309; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid310_In0 <= "" & bh4_w5_50 & bh4_w5_47 & bh4_w5_45 & bh4_w5_43 & bh4_w5_48 & bh4_w5_49;
   bh4_w5_54 <= Compressor_6_3_F125_uid69_bh4_uid310_Out0(0);
   bh4_w6_49 <= Compressor_6_3_F125_uid69_bh4_uid310_Out0(1);
   bh4_w7_44 <= Compressor_6_3_F125_uid69_bh4_uid310_Out0(2);
   Compressor_6_3_F125_uid69_uid310: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid310_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid310_Out0_copy311);
   Compressor_6_3_F125_uid69_bh4_uid310_Out0 <= Compressor_6_3_F125_uid69_bh4_uid310_Out0_copy311; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid312_In0 <= "" & bh4_w5_34 & bh4_w5_44 & bh4_w5_46;
   Compressor_23_3_F125_uid193_bh4_uid312_In1 <= "" & bh4_w6_47 & bh4_w6_43;
   bh4_w5_55 <= Compressor_23_3_F125_uid193_bh4_uid312_Out0(0);
   bh4_w6_50 <= Compressor_23_3_F125_uid193_bh4_uid312_Out0(1);
   bh4_w7_45 <= Compressor_23_3_F125_uid193_bh4_uid312_Out0(2);
   Compressor_23_3_F125_uid193_uid312: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid312_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid312_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid312_Out0_copy313);
   Compressor_23_3_F125_uid193_bh4_uid312_Out0 <= Compressor_23_3_F125_uid193_bh4_uid312_Out0_copy313; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid314_In0 <= "" & bh4_w6_41 & bh4_w6_45 & bh4_w6_46 & bh4_w6_40 & bh4_w6_42 & bh4_w6_44;
   bh4_w6_51 <= Compressor_6_3_F125_uid69_bh4_uid314_Out0(0);
   bh4_w7_46 <= Compressor_6_3_F125_uid69_bh4_uid314_Out0(1);
   bh4_w8_40 <= Compressor_6_3_F125_uid69_bh4_uid314_Out0(2);
   Compressor_6_3_F125_uid69_uid314: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid314_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid314_Out0_copy315);
   Compressor_6_3_F125_uid69_bh4_uid314_Out0 <= Compressor_6_3_F125_uid69_bh4_uid314_Out0_copy315; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid316_In0 <= "" & bh4_w7_41 & bh4_w7_39 & bh4_w7_38 & bh4_w7_37 & bh4_w7_42 & "0";
   bh4_w7_47 <= Compressor_6_3_F125_uid69_bh4_uid316_Out0(0);
   bh4_w8_41 <= Compressor_6_3_F125_uid69_bh4_uid316_Out0(1);
   bh4_w9_37 <= Compressor_6_3_F125_uid69_bh4_uid316_Out0(2);
   Compressor_6_3_F125_uid69_uid316: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid316_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid316_Out0_copy317);
   Compressor_6_3_F125_uid69_bh4_uid316_Out0 <= Compressor_6_3_F125_uid69_bh4_uid316_Out0_copy317; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid318_In0 <= "" & bh4_w7_43 & bh4_w7_28 & bh4_w7_40;
   bh4_w7_48 <= Compressor_3_2_F125_uid223_bh4_uid318_Out0(0);
   bh4_w8_42 <= Compressor_3_2_F125_uid223_bh4_uid318_Out0(1);
   Compressor_3_2_F125_uid223_uid318: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid318_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid318_Out0_copy319);
   Compressor_3_2_F125_uid223_bh4_uid318_Out0 <= Compressor_3_2_F125_uid223_bh4_uid318_Out0_copy319; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid320_In0 <= "" & bh4_w8_37 & bh4_w8_36 & bh4_w8_35 & bh4_w8_34 & bh4_w8_38 & bh4_w8_39;
   bh4_w8_43 <= Compressor_6_3_F125_uid69_bh4_uid320_Out0(0);
   bh4_w9_38 <= Compressor_6_3_F125_uid69_bh4_uid320_Out0(1);
   bh4_w10_34 <= Compressor_6_3_F125_uid69_bh4_uid320_Out0(2);
   Compressor_6_3_F125_uid69_uid320: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid320_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid320_Out0_copy321);
   Compressor_6_3_F125_uid69_bh4_uid320_Out0 <= Compressor_6_3_F125_uid69_bh4_uid320_Out0_copy321; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid322_In0 <= "" & bh4_w9_34 & bh4_w9_33 & bh4_w9_32 & bh4_w9_31 & bh4_w9_35 & bh4_w9_36;
   bh4_w9_39 <= Compressor_6_3_F125_uid69_bh4_uid322_Out0(0);
   bh4_w10_35 <= Compressor_6_3_F125_uid69_bh4_uid322_Out0(1);
   bh4_w11_31 <= Compressor_6_3_F125_uid69_bh4_uid322_Out0(2);
   Compressor_6_3_F125_uid69_uid322: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid322_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid322_Out0_copy323);
   Compressor_6_3_F125_uid69_bh4_uid322_Out0 <= Compressor_6_3_F125_uid69_bh4_uid322_Out0_copy323; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid324_In0 <= "" & bh4_w10_33 & bh4_w10_32 & bh4_w10_31 & bh4_w10_30 & bh4_w10_29 & bh4_w10_28;
   bh4_w10_36 <= Compressor_6_3_F125_uid69_bh4_uid324_Out0(0);
   bh4_w11_32 <= Compressor_6_3_F125_uid69_bh4_uid324_Out0(1);
   bh4_w12_28 <= Compressor_6_3_F125_uid69_bh4_uid324_Out0(2);
   Compressor_6_3_F125_uid69_uid324: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid324_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid324_Out0_copy325);
   Compressor_6_3_F125_uid69_bh4_uid324_Out0 <= Compressor_6_3_F125_uid69_bh4_uid324_Out0_copy325; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid326_In0 <= "" & bh4_w11_30 & bh4_w11_29 & bh4_w11_28 & bh4_w11_27 & bh4_w11_26 & bh4_w11_25;
   bh4_w11_33 <= Compressor_6_3_F125_uid69_bh4_uid326_Out0(0);
   bh4_w12_29 <= Compressor_6_3_F125_uid69_bh4_uid326_Out0(1);
   bh4_w13_23 <= Compressor_6_3_F125_uid69_bh4_uid326_Out0(2);
   Compressor_6_3_F125_uid69_uid326: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid326_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid326_Out0_copy327);
   Compressor_6_3_F125_uid69_bh4_uid326_Out0 <= Compressor_6_3_F125_uid69_bh4_uid326_Out0_copy327; -- output copy to hold a pipeline register if needed


   Compressor_6_3_F125_uid69_bh4_uid328_In0 <= "" & bh4_w12_27 & bh4_w12_26 & bh4_w12_25 & bh4_w12_24 & bh4_w12_23 & bh4_w12_22;
   bh4_w12_30 <= Compressor_6_3_F125_uid69_bh4_uid328_Out0(0);
   bh4_w13_24 <= Compressor_6_3_F125_uid69_bh4_uid328_Out0(1);
   bh4_w14_19 <= Compressor_6_3_F125_uid69_bh4_uid328_Out0(2);
   Compressor_6_3_F125_uid69_uid328: Compressor_6_3_F125_uid69
      port map ( X0 => Compressor_6_3_F125_uid69_bh4_uid328_In0,
                 R => Compressor_6_3_F125_uid69_bh4_uid328_Out0_copy329);
   Compressor_6_3_F125_uid69_bh4_uid328_Out0 <= Compressor_6_3_F125_uid69_bh4_uid328_Out0_copy329; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid330_In0 <= "" & bh4_w13_22 & bh4_w13_21 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid330_In1 <= "" & bh4_w14_18;
   bh4_w13_25 <= Compressor_14_3_F125_uid79_bh4_uid330_Out0(0);
   bh4_w14_20 <= Compressor_14_3_F125_uid79_bh4_uid330_Out0(1);
   bh4_w15_16 <= Compressor_14_3_F125_uid79_bh4_uid330_Out0(2);
   Compressor_14_3_F125_uid79_uid330: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid330_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid330_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid330_Out0_copy331);
   Compressor_14_3_F125_uid79_bh4_uid330_Out0 <= Compressor_14_3_F125_uid79_bh4_uid330_Out0_copy331; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid332_In0 <= "" & bh4_w13_20 & bh4_w13_19 & bh4_w13_18;
   Compressor_23_3_F125_uid193_bh4_uid332_In1 <= "" & bh4_w14_17 & bh4_w14_16;
   bh4_w13_26 <= Compressor_23_3_F125_uid193_bh4_uid332_Out0(0);
   bh4_w14_21 <= Compressor_23_3_F125_uid193_bh4_uid332_Out0(1);
   bh4_w15_17 <= Compressor_23_3_F125_uid193_bh4_uid332_Out0(2);
   Compressor_23_3_F125_uid193_uid332: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid332_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid332_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid332_Out0_copy333);
   Compressor_23_3_F125_uid193_bh4_uid332_Out0 <= Compressor_23_3_F125_uid193_bh4_uid332_Out0_copy333; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid334_In0 <= "" & bh4_w15_15 & bh4_w15_14 & bh4_w15_13;
   Compressor_23_3_F125_uid193_bh4_uid334_In1 <= "" & bh4_w16_12 & bh4_w16_11;
   bh4_w15_18 <= Compressor_23_3_F125_uid193_bh4_uid334_Out0(0);
   bh4_w16_13 <= Compressor_23_3_F125_uid193_bh4_uid334_Out0(1);
   bh4_w17_11 <= Compressor_23_3_F125_uid193_bh4_uid334_Out0(2);
   Compressor_23_3_F125_uid193_uid334: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid334_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid334_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid334_Out0_copy335);
   Compressor_23_3_F125_uid193_bh4_uid334_Out0 <= Compressor_23_3_F125_uid193_bh4_uid334_Out0_copy335; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid336_In0 <= "" & bh4_w17_10 & bh4_w17_9 & bh4_w17_8;
   Compressor_23_3_F125_uid193_bh4_uid336_In1 <= "" & bh4_w18_7 & bh4_w18_6;
   bh4_w17_12 <= Compressor_23_3_F125_uid193_bh4_uid336_Out0(0);
   bh4_w18_8 <= Compressor_23_3_F125_uid193_bh4_uid336_Out0(1);
   bh4_w19_6 <= Compressor_23_3_F125_uid193_bh4_uid336_Out0(2);
   Compressor_23_3_F125_uid193_uid336: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid336_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid336_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid336_Out0_copy337);
   Compressor_23_3_F125_uid193_bh4_uid336_Out0 <= Compressor_23_3_F125_uid193_bh4_uid336_Out0_copy337; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid338_In0 <= "" & bh4_w19_5 & bh4_w19_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid338_In1 <= "" & bh4_w20_4;
   bh4_w19_7 <= Compressor_14_3_F125_uid79_bh4_uid338_Out0(0);
   bh4_w20_5 <= Compressor_14_3_F125_uid79_bh4_uid338_Out0(1);
   bh4_w21_4 <= Compressor_14_3_F125_uid79_bh4_uid338_Out0(2);
   Compressor_14_3_F125_uid79_uid338: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid338_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid338_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid338_Out0_copy339);
   Compressor_14_3_F125_uid79_bh4_uid338_Out0 <= Compressor_14_3_F125_uid79_bh4_uid338_Out0_copy339; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid340_In0 <= "" & bh4_w21_3 & bh4_w21_2 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid340_In1 <= "" & bh4_w22_4;
   bh4_w21_5 <= Compressor_14_3_F125_uid79_bh4_uid340_Out0(0);
   bh4_w22_5 <= Compressor_14_3_F125_uid79_bh4_uid340_Out0(1);
   bh4_w23_4 <= Compressor_14_3_F125_uid79_bh4_uid340_Out0(2);
   Compressor_14_3_F125_uid79_uid340: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid340_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid340_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid340_Out0_copy341);
   Compressor_14_3_F125_uid79_bh4_uid340_Out0 <= Compressor_14_3_F125_uid79_bh4_uid340_Out0_copy341; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid342_In0 <= "" & bh4_w24_5 & bh4_w24_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid342_In1 <= "" & bh4_w25_3;
   bh4_w24_6 <= Compressor_14_3_F125_uid79_bh4_uid342_Out0(0);
   bh4_w25_4 <= Compressor_14_3_F125_uid79_bh4_uid342_Out0(1);
   bh4_w26_6 <= Compressor_14_3_F125_uid79_bh4_uid342_Out0(2);
   Compressor_14_3_F125_uid79_uid342: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid342_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid342_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid342_Out0_copy343);
   Compressor_14_3_F125_uid79_bh4_uid342_Out0 <= Compressor_14_3_F125_uid79_bh4_uid342_Out0_copy343; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid344_In0 <= "" & bh4_w26_5 & bh4_w26_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid344_In1 <= "" & bh4_w27_3;
   bh4_w26_7 <= Compressor_14_3_F125_uid79_bh4_uid344_Out0(0);
   bh4_w27_4 <= Compressor_14_3_F125_uid79_bh4_uid344_Out0(1);
   bh4_w28_6 <= Compressor_14_3_F125_uid79_bh4_uid344_Out0(2);
   Compressor_14_3_F125_uid79_uid344: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid344_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid344_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid344_Out0_copy345);
   Compressor_14_3_F125_uid79_bh4_uid344_Out0 <= Compressor_14_3_F125_uid79_bh4_uid344_Out0_copy345; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid346_In0 <= "" & bh4_w28_5 & bh4_w28_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid346_In1 <= "" & bh4_w29_3;
   bh4_w28_7 <= Compressor_14_3_F125_uid79_bh4_uid346_Out0(0);
   bh4_w29_4 <= Compressor_14_3_F125_uid79_bh4_uid346_Out0(1);
   bh4_w30_6 <= Compressor_14_3_F125_uid79_bh4_uid346_Out0(2);
   Compressor_14_3_F125_uid79_uid346: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid346_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid346_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid346_Out0_copy347);
   Compressor_14_3_F125_uid79_bh4_uid346_Out0 <= Compressor_14_3_F125_uid79_bh4_uid346_Out0_copy347; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid348_In0 <= "" & bh4_w30_5 & bh4_w30_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid348_In1 <= "" & bh4_w31_3;
   bh4_w30_7 <= Compressor_14_3_F125_uid79_bh4_uid348_Out0(0);
   bh4_w31_4 <= Compressor_14_3_F125_uid79_bh4_uid348_Out0(1);
   bh4_w32_6 <= Compressor_14_3_F125_uid79_bh4_uid348_Out0(2);
   Compressor_14_3_F125_uid79_uid348: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid348_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid348_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid348_Out0_copy349);
   Compressor_14_3_F125_uid79_bh4_uid348_Out0 <= Compressor_14_3_F125_uid79_bh4_uid348_Out0_copy349; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid350_In0 <= "" & bh4_w32_5 & bh4_w32_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid350_In1 <= "" & bh4_w33_3;
   bh4_w32_7 <= Compressor_14_3_F125_uid79_bh4_uid350_Out0(0);
   bh4_w33_4 <= Compressor_14_3_F125_uid79_bh4_uid350_Out0(1);
   bh4_w34_6 <= Compressor_14_3_F125_uid79_bh4_uid350_Out0(2);
   Compressor_14_3_F125_uid79_uid350: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid350_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid350_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid350_Out0_copy351);
   Compressor_14_3_F125_uid79_bh4_uid350_Out0 <= Compressor_14_3_F125_uid79_bh4_uid350_Out0_copy351; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid352_In0 <= "" & bh4_w34_5 & bh4_w34_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid352_In1 <= "" & bh4_w35_3;
   bh4_w34_7 <= Compressor_14_3_F125_uid79_bh4_uid352_Out0(0);
   bh4_w35_4 <= Compressor_14_3_F125_uid79_bh4_uid352_Out0(1);
   bh4_w36_4 <= Compressor_14_3_F125_uid79_bh4_uid352_Out0(2);
   Compressor_14_3_F125_uid79_uid352: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid352_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid352_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid352_Out0_copy353);
   Compressor_14_3_F125_uid79_bh4_uid352_Out0 <= Compressor_14_3_F125_uid79_bh4_uid352_Out0_copy353; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid354_In0 <= "" & bh4_w36_3 & bh4_w36_2 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid354_In1 <= "" & bh4_w37_1;
   bh4_w36_5 <= Compressor_14_3_F125_uid79_bh4_uid354_Out0(0);
   bh4_w37_2 <= Compressor_14_3_F125_uid79_bh4_uid354_Out0(1);
   bh4_w38_2 <= Compressor_14_3_F125_uid79_bh4_uid354_Out0(2);
   Compressor_14_3_F125_uid79_uid354: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid354_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid354_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid354_Out0_copy355);
   Compressor_14_3_F125_uid79_bh4_uid354_Out0 <= Compressor_14_3_F125_uid79_bh4_uid354_Out0_copy355; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid356_In0 <= "" & bh4_w38_0 & bh4_w38_1 & "0";
   bh4_w38_3 <= Compressor_3_2_F125_uid223_bh4_uid356_Out0(0);
   bh4_w39_0 <= Compressor_3_2_F125_uid223_bh4_uid356_Out0(1);
   Compressor_3_2_F125_uid223_uid356: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid356_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid356_Out0_copy357);
   Compressor_3_2_F125_uid223_bh4_uid356_Out0 <= Compressor_3_2_F125_uid223_bh4_uid356_Out0_copy357; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid358_In0 <= "" & bh4_w1_44 & "0" & "0";
   Compressor_23_3_F125_uid193_bh4_uid358_In1 <= "" & bh4_w2_53 & bh4_w2_52;
   bh4_w1_45 <= Compressor_23_3_F125_uid193_bh4_uid358_Out0(0);
   bh4_w2_54 <= Compressor_23_3_F125_uid193_bh4_uid358_Out0(1);
   bh4_w3_57 <= Compressor_23_3_F125_uid193_bh4_uid358_Out0(2);
   Compressor_23_3_F125_uid193_uid358: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid358_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid358_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid358_Out0_copy359);
   Compressor_23_3_F125_uid193_bh4_uid358_Out0 <= Compressor_23_3_F125_uid193_bh4_uid358_Out0_copy359; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid360_In0 <= "" & bh4_w3_56 & bh4_w3_55 & bh4_w3_54;
   bh4_w3_58 <= Compressor_3_2_F125_uid223_bh4_uid360_Out0(0);
   bh4_w4_58 <= Compressor_3_2_F125_uid223_bh4_uid360_Out0(1);
   Compressor_3_2_F125_uid223_uid360: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid360_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid360_Out0_copy361);
   Compressor_3_2_F125_uid223_bh4_uid360_Out0 <= Compressor_3_2_F125_uid223_bh4_uid360_Out0_copy361; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid362_In0 <= "" & bh4_w4_57 & bh4_w4_56 & bh4_w4_55 & bh4_w4_54;
   Compressor_14_3_F125_uid79_bh4_uid362_In1 <= "" & bh4_w5_55;
   bh4_w4_59 <= Compressor_14_3_F125_uid79_bh4_uid362_Out0(0);
   bh4_w5_56 <= Compressor_14_3_F125_uid79_bh4_uid362_Out0(1);
   bh4_w6_52 <= Compressor_14_3_F125_uid79_bh4_uid362_Out0(2);
   Compressor_14_3_F125_uid79_uid362: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid362_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid362_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid362_Out0_copy363);
   Compressor_14_3_F125_uid79_bh4_uid362_Out0 <= Compressor_14_3_F125_uid79_bh4_uid362_Out0_copy363; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid364_In0 <= "" & bh4_w5_54 & bh4_w5_53 & bh4_w5_52 & bh4_w5_51;
   Compressor_14_3_F125_uid79_bh4_uid364_In1 <= "" & bh4_w6_51;
   bh4_w5_57 <= Compressor_14_3_F125_uid79_bh4_uid364_Out0(0);
   bh4_w6_53 <= Compressor_14_3_F125_uid79_bh4_uid364_Out0(1);
   bh4_w7_49 <= Compressor_14_3_F125_uid79_bh4_uid364_Out0(2);
   Compressor_14_3_F125_uid79_uid364: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid364_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid364_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid364_Out0_copy365);
   Compressor_14_3_F125_uid79_bh4_uid364_Out0 <= Compressor_14_3_F125_uid79_bh4_uid364_Out0_copy365; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid366_In0 <= "" & bh4_w6_50 & bh4_w6_49 & bh4_w6_48;
   bh4_w6_54 <= Compressor_3_2_F125_uid223_bh4_uid366_Out0(0);
   bh4_w7_50 <= Compressor_3_2_F125_uid223_bh4_uid366_Out0(1);
   Compressor_3_2_F125_uid223_uid366: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid366_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid366_Out0_copy367);
   Compressor_3_2_F125_uid223_bh4_uid366_Out0 <= Compressor_3_2_F125_uid223_bh4_uid366_Out0_copy367; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid368_In0 <= "" & bh4_w7_48 & bh4_w7_47 & bh4_w7_46 & bh4_w7_45;
   Compressor_14_3_F125_uid79_bh4_uid368_In1 <= "" & bh4_w8_43;
   bh4_w7_51 <= Compressor_14_3_F125_uid79_bh4_uid368_Out0(0);
   bh4_w8_44 <= Compressor_14_3_F125_uid79_bh4_uid368_Out0(1);
   bh4_w9_40 <= Compressor_14_3_F125_uid79_bh4_uid368_Out0(2);
   Compressor_14_3_F125_uid79_uid368: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid368_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid368_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid368_Out0_copy369);
   Compressor_14_3_F125_uid79_bh4_uid368_Out0 <= Compressor_14_3_F125_uid79_bh4_uid368_Out0_copy369; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid370_In0 <= "" & bh4_w8_42 & bh4_w8_41 & bh4_w8_40;
   Compressor_23_3_F125_uid193_bh4_uid370_In1 <= "" & bh4_w9_39 & bh4_w9_38;
   bh4_w8_45 <= Compressor_23_3_F125_uid193_bh4_uid370_Out0(0);
   bh4_w9_41 <= Compressor_23_3_F125_uid193_bh4_uid370_Out0(1);
   bh4_w10_37 <= Compressor_23_3_F125_uid193_bh4_uid370_Out0(2);
   Compressor_23_3_F125_uid193_uid370: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid370_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid370_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid370_Out0_copy371);
   Compressor_23_3_F125_uid193_bh4_uid370_Out0 <= Compressor_23_3_F125_uid193_bh4_uid370_Out0_copy371; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid372_In0 <= "" & bh4_w10_36 & bh4_w10_35 & bh4_w10_34;
   Compressor_23_3_F125_uid193_bh4_uid372_In1 <= "" & bh4_w11_33 & bh4_w11_32;
   bh4_w10_38 <= Compressor_23_3_F125_uid193_bh4_uid372_Out0(0);
   bh4_w11_34 <= Compressor_23_3_F125_uid193_bh4_uid372_Out0(1);
   bh4_w12_31 <= Compressor_23_3_F125_uid193_bh4_uid372_Out0(2);
   Compressor_23_3_F125_uid193_uid372: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid372_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid372_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid372_Out0_copy373);
   Compressor_23_3_F125_uid193_bh4_uid372_Out0 <= Compressor_23_3_F125_uid193_bh4_uid372_Out0_copy373; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid374_In0 <= "" & bh4_w12_30 & bh4_w12_29 & bh4_w12_28;
   bh4_w12_32 <= Compressor_3_2_F125_uid223_bh4_uid374_Out0(0);
   bh4_w13_27 <= Compressor_3_2_F125_uid223_bh4_uid374_Out0(1);
   Compressor_3_2_F125_uid223_uid374: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid374_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid374_Out0_copy375);
   Compressor_3_2_F125_uid223_bh4_uid374_Out0 <= Compressor_3_2_F125_uid223_bh4_uid374_Out0_copy375; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid376_In0 <= "" & bh4_w13_26 & bh4_w13_25 & bh4_w13_24 & bh4_w13_23;
   Compressor_14_3_F125_uid79_bh4_uid376_In1 <= "" & "0";
   bh4_w13_28 <= Compressor_14_3_F125_uid79_bh4_uid376_Out0(0);
   bh4_w14_22 <= Compressor_14_3_F125_uid79_bh4_uid376_Out0(1);
   bh4_w15_19 <= Compressor_14_3_F125_uid79_bh4_uid376_Out0(2);
   Compressor_14_3_F125_uid79_uid376: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid376_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid376_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid376_Out0_copy377);
   Compressor_14_3_F125_uid79_bh4_uid376_Out0 <= Compressor_14_3_F125_uid79_bh4_uid376_Out0_copy377; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid378_In0 <= "" & bh4_w14_21 & bh4_w14_20 & bh4_w14_19;
   bh4_w14_23 <= Compressor_3_2_F125_uid223_bh4_uid378_Out0(0);
   bh4_w15_20 <= Compressor_3_2_F125_uid223_bh4_uid378_Out0(1);
   Compressor_3_2_F125_uid223_uid378: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid378_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid378_Out0_copy379);
   Compressor_3_2_F125_uid223_bh4_uid378_Out0 <= Compressor_3_2_F125_uid223_bh4_uid378_Out0_copy379; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid380_In0 <= "" & bh4_w15_18 & bh4_w15_17 & bh4_w15_16;
   Compressor_23_3_F125_uid193_bh4_uid380_In1 <= "" & bh4_w16_13 & bh4_w16_10;
   bh4_w15_21 <= Compressor_23_3_F125_uid193_bh4_uid380_Out0(0);
   bh4_w16_14 <= Compressor_23_3_F125_uid193_bh4_uid380_Out0(1);
   bh4_w17_13 <= Compressor_23_3_F125_uid193_bh4_uid380_Out0(2);
   Compressor_23_3_F125_uid193_uid380: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid380_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid380_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid380_Out0_copy381);
   Compressor_23_3_F125_uid193_bh4_uid380_Out0 <= Compressor_23_3_F125_uid193_bh4_uid380_Out0_copy381; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid382_In0 <= "" & bh4_w17_12 & bh4_w17_11 & "0";
   Compressor_23_3_F125_uid193_bh4_uid382_In1 <= "" & bh4_w18_8 & bh4_w18_3;
   bh4_w17_14 <= Compressor_23_3_F125_uid193_bh4_uid382_Out0(0);
   bh4_w18_9 <= Compressor_23_3_F125_uid193_bh4_uid382_Out0(1);
   bh4_w19_8 <= Compressor_23_3_F125_uid193_bh4_uid382_Out0(2);
   Compressor_23_3_F125_uid193_uid382: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid382_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid382_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid382_Out0_copy383);
   Compressor_23_3_F125_uid193_bh4_uid382_Out0 <= Compressor_23_3_F125_uid193_bh4_uid382_Out0_copy383; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid384_In0 <= "" & bh4_w19_7 & bh4_w19_6 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid384_In1 <= "" & bh4_w20_5;
   bh4_w19_9 <= Compressor_14_3_F125_uid79_bh4_uid384_Out0(0);
   bh4_w20_6 <= Compressor_14_3_F125_uid79_bh4_uid384_Out0(1);
   bh4_w21_6 <= Compressor_14_3_F125_uid79_bh4_uid384_Out0(2);
   Compressor_14_3_F125_uid79_uid384: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid384_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid384_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid384_Out0_copy385);
   Compressor_14_3_F125_uid79_bh4_uid384_Out0 <= Compressor_14_3_F125_uid79_bh4_uid384_Out0_copy385; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid386_In0 <= "" & bh4_w21_5 & bh4_w21_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid386_In1 <= "" & bh4_w22_5;
   bh4_w21_7 <= Compressor_14_3_F125_uid79_bh4_uid386_Out0(0);
   bh4_w22_6 <= Compressor_14_3_F125_uid79_bh4_uid386_Out0(1);
   bh4_w23_5 <= Compressor_14_3_F125_uid79_bh4_uid386_Out0(2);
   Compressor_14_3_F125_uid79_uid386: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid386_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid386_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid386_Out0_copy387);
   Compressor_14_3_F125_uid79_bh4_uid386_Out0 <= Compressor_14_3_F125_uid79_bh4_uid386_Out0_copy387; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid388_In0 <= "" & bh4_w23_4 & bh4_w23_3 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid388_In1 <= "" & bh4_w24_6;
   bh4_w23_6 <= Compressor_14_3_F125_uid79_bh4_uid388_Out0(0);
   bh4_w24_7 <= Compressor_14_3_F125_uid79_bh4_uid388_Out0(1);
   bh4_w25_5 <= Compressor_14_3_F125_uid79_bh4_uid388_Out0(2);
   Compressor_14_3_F125_uid79_uid388: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid388_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid388_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid388_Out0_copy389);
   Compressor_14_3_F125_uid79_bh4_uid388_Out0 <= Compressor_14_3_F125_uid79_bh4_uid388_Out0_copy389; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid390_In0 <= "" & bh4_w26_7 & bh4_w26_6 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid390_In1 <= "" & bh4_w27_4;
   bh4_w26_8 <= Compressor_14_3_F125_uid79_bh4_uid390_Out0(0);
   bh4_w27_5 <= Compressor_14_3_F125_uid79_bh4_uid390_Out0(1);
   bh4_w28_8 <= Compressor_14_3_F125_uid79_bh4_uid390_Out0(2);
   Compressor_14_3_F125_uid79_uid390: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid390_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid390_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid390_Out0_copy391);
   Compressor_14_3_F125_uid79_bh4_uid390_Out0 <= Compressor_14_3_F125_uid79_bh4_uid390_Out0_copy391; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid392_In0 <= "" & bh4_w28_7 & bh4_w28_6 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid392_In1 <= "" & bh4_w29_4;
   bh4_w28_9 <= Compressor_14_3_F125_uid79_bh4_uid392_Out0(0);
   bh4_w29_5 <= Compressor_14_3_F125_uid79_bh4_uid392_Out0(1);
   bh4_w30_8 <= Compressor_14_3_F125_uid79_bh4_uid392_Out0(2);
   Compressor_14_3_F125_uid79_uid392: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid392_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid392_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid392_Out0_copy393);
   Compressor_14_3_F125_uid79_bh4_uid392_Out0 <= Compressor_14_3_F125_uid79_bh4_uid392_Out0_copy393; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid394_In0 <= "" & bh4_w30_7 & bh4_w30_6 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid394_In1 <= "" & bh4_w31_4;
   bh4_w30_9 <= Compressor_14_3_F125_uid79_bh4_uid394_Out0(0);
   bh4_w31_5 <= Compressor_14_3_F125_uid79_bh4_uid394_Out0(1);
   bh4_w32_8 <= Compressor_14_3_F125_uid79_bh4_uid394_Out0(2);
   Compressor_14_3_F125_uid79_uid394: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid394_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid394_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid394_Out0_copy395);
   Compressor_14_3_F125_uid79_bh4_uid394_Out0 <= Compressor_14_3_F125_uid79_bh4_uid394_Out0_copy395; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid396_In0 <= "" & bh4_w32_7 & bh4_w32_6 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid396_In1 <= "" & bh4_w33_4;
   bh4_w32_9 <= Compressor_14_3_F125_uid79_bh4_uid396_Out0(0);
   bh4_w33_5 <= Compressor_14_3_F125_uid79_bh4_uid396_Out0(1);
   bh4_w34_8 <= Compressor_14_3_F125_uid79_bh4_uid396_Out0(2);
   Compressor_14_3_F125_uid79_uid396: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid396_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid396_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid396_Out0_copy397);
   Compressor_14_3_F125_uid79_bh4_uid396_Out0 <= Compressor_14_3_F125_uid79_bh4_uid396_Out0_copy397; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid398_In0 <= "" & bh4_w34_7 & bh4_w34_6 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid398_In1 <= "" & bh4_w35_4;
   bh4_w34_9 <= Compressor_14_3_F125_uid79_bh4_uid398_Out0(0);
   bh4_w35_5 <= Compressor_14_3_F125_uid79_bh4_uid398_Out0(1);
   bh4_w36_6 <= Compressor_14_3_F125_uid79_bh4_uid398_Out0(2);
   Compressor_14_3_F125_uid79_uid398: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid398_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid398_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid398_Out0_copy399);
   Compressor_14_3_F125_uid79_bh4_uid398_Out0 <= Compressor_14_3_F125_uid79_bh4_uid398_Out0_copy399; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid400_In0 <= "" & bh4_w36_5 & bh4_w36_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid400_In1 <= "" & bh4_w37_2;
   bh4_w36_7 <= Compressor_14_3_F125_uid79_bh4_uid400_Out0(0);
   bh4_w37_3 <= Compressor_14_3_F125_uid79_bh4_uid400_Out0(1);
   bh4_w38_4 <= Compressor_14_3_F125_uid79_bh4_uid400_Out0(2);
   Compressor_14_3_F125_uid79_uid400: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid400_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid400_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid400_Out0_copy401);
   Compressor_14_3_F125_uid79_bh4_uid400_Out0 <= Compressor_14_3_F125_uid79_bh4_uid400_Out0_copy401; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid402_In0 <= "" & bh4_w38_3 & bh4_w38_2 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid402_In1 <= "" & bh4_w39_0;
   bh4_w38_5 <= Compressor_14_3_F125_uid79_bh4_uid402_Out0(0);
   bh4_w39_1 <= Compressor_14_3_F125_uid79_bh4_uid402_Out0(1);
   bh4_w40_0 <= Compressor_14_3_F125_uid79_bh4_uid402_Out0(2);
   Compressor_14_3_F125_uid79_uid402: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid402_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid402_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid402_Out0_copy403);
   Compressor_14_3_F125_uid79_bh4_uid402_Out0 <= Compressor_14_3_F125_uid79_bh4_uid402_Out0_copy403; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid404_In0 <= "" & bh4_w3_58 & bh4_w3_57 & "0";
   Compressor_23_3_F125_uid193_bh4_uid404_In1 <= "" & bh4_w4_59 & bh4_w4_58;
   bh4_w3_59 <= Compressor_23_3_F125_uid193_bh4_uid404_Out0(0);
   bh4_w4_60 <= Compressor_23_3_F125_uid193_bh4_uid404_Out0(1);
   bh4_w5_58 <= Compressor_23_3_F125_uid193_bh4_uid404_Out0(2);
   Compressor_23_3_F125_uid193_uid404: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid404_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid404_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid404_Out0_copy405);
   Compressor_23_3_F125_uid193_bh4_uid404_Out0 <= Compressor_23_3_F125_uid193_bh4_uid404_Out0_copy405; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid406_In0 <= "" & bh4_w5_57 & bh4_w5_56 & "0";
   bh4_w5_59 <= Compressor_3_2_F125_uid223_bh4_uid406_Out0(0);
   bh4_w6_55 <= Compressor_3_2_F125_uid223_bh4_uid406_Out0(1);
   Compressor_3_2_F125_uid223_uid406: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid406_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid406_Out0_copy407);
   Compressor_3_2_F125_uid223_bh4_uid406_Out0 <= Compressor_3_2_F125_uid223_bh4_uid406_Out0_copy407; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid408_In0 <= "" & bh4_w6_54 & bh4_w6_53 & bh4_w6_52;
   bh4_w6_56 <= Compressor_3_2_F125_uid223_bh4_uid408_Out0(0);
   bh4_w7_52 <= Compressor_3_2_F125_uid223_bh4_uid408_Out0(1);
   Compressor_3_2_F125_uid223_uid408: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid408_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid408_Out0_copy409);
   Compressor_3_2_F125_uid223_bh4_uid408_Out0 <= Compressor_3_2_F125_uid223_bh4_uid408_Out0_copy409; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid410_In0 <= "" & bh4_w7_51 & bh4_w7_50 & bh4_w7_49 & bh4_w7_44;
   Compressor_14_3_F125_uid79_bh4_uid410_In1 <= "" & bh4_w8_45;
   bh4_w7_53 <= Compressor_14_3_F125_uid79_bh4_uid410_Out0(0);
   bh4_w8_46 <= Compressor_14_3_F125_uid79_bh4_uid410_Out0(1);
   bh4_w9_42 <= Compressor_14_3_F125_uid79_bh4_uid410_Out0(2);
   Compressor_14_3_F125_uid79_uid410: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid410_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid410_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid410_Out0_copy411);
   Compressor_14_3_F125_uid79_bh4_uid410_Out0 <= Compressor_14_3_F125_uid79_bh4_uid410_Out0_copy411; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid412_In0 <= "" & bh4_w9_41 & bh4_w9_40 & bh4_w9_37;
   Compressor_23_3_F125_uid193_bh4_uid412_In1 <= "" & bh4_w10_38 & bh4_w10_37;
   bh4_w9_43 <= Compressor_23_3_F125_uid193_bh4_uid412_Out0(0);
   bh4_w10_39 <= Compressor_23_3_F125_uid193_bh4_uid412_Out0(1);
   bh4_w11_35 <= Compressor_23_3_F125_uid193_bh4_uid412_Out0(2);
   Compressor_23_3_F125_uid193_uid412: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid412_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid412_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid412_Out0_copy413);
   Compressor_23_3_F125_uid193_bh4_uid412_Out0 <= Compressor_23_3_F125_uid193_bh4_uid412_Out0_copy413; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid414_In0 <= "" & bh4_w11_34 & bh4_w11_31 & "0";
   Compressor_23_3_F125_uid193_bh4_uid414_In1 <= "" & bh4_w12_32 & bh4_w12_31;
   bh4_w11_36 <= Compressor_23_3_F125_uid193_bh4_uid414_Out0(0);
   bh4_w12_33 <= Compressor_23_3_F125_uid193_bh4_uid414_Out0(1);
   bh4_w13_29 <= Compressor_23_3_F125_uid193_bh4_uid414_Out0(2);
   Compressor_23_3_F125_uid193_uid414: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid414_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid414_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid414_Out0_copy415);
   Compressor_23_3_F125_uid193_bh4_uid414_Out0 <= Compressor_23_3_F125_uid193_bh4_uid414_Out0_copy415; -- output copy to hold a pipeline register if needed


   Compressor_23_3_F125_uid193_bh4_uid416_In0 <= "" & bh4_w13_28 & bh4_w13_27 & "0";
   Compressor_23_3_F125_uid193_bh4_uid416_In1 <= "" & bh4_w14_23 & bh4_w14_22;
   bh4_w13_30 <= Compressor_23_3_F125_uid193_bh4_uid416_Out0(0);
   bh4_w14_24 <= Compressor_23_3_F125_uid193_bh4_uid416_Out0(1);
   bh4_w15_22 <= Compressor_23_3_F125_uid193_bh4_uid416_Out0(2);
   Compressor_23_3_F125_uid193_uid416: Compressor_23_3_F125_uid193
      port map ( X0 => Compressor_23_3_F125_uid193_bh4_uid416_In0,
                 X1 => Compressor_23_3_F125_uid193_bh4_uid416_In1,
                 R => Compressor_23_3_F125_uid193_bh4_uid416_Out0_copy417);
   Compressor_23_3_F125_uid193_bh4_uid416_Out0 <= Compressor_23_3_F125_uid193_bh4_uid416_Out0_copy417; -- output copy to hold a pipeline register if needed


   Compressor_3_2_F125_uid223_bh4_uid418_In0 <= "" & bh4_w15_21 & bh4_w15_20 & bh4_w15_19;
   bh4_w15_23 <= Compressor_3_2_F125_uid223_bh4_uid418_Out0(0);
   bh4_w16_15 <= Compressor_3_2_F125_uid223_bh4_uid418_Out0(1);
   Compressor_3_2_F125_uid223_uid418: Compressor_3_2_F125_uid223
      port map ( X0 => Compressor_3_2_F125_uid223_bh4_uid418_In0,
                 R => Compressor_3_2_F125_uid223_bh4_uid418_Out0_copy419);
   Compressor_3_2_F125_uid223_bh4_uid418_Out0 <= Compressor_3_2_F125_uid223_bh4_uid418_Out0_copy419; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid420_In0 <= "" & bh4_w17_14 & bh4_w17_13 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid420_In1 <= "" & bh4_w18_9;
   bh4_w17_15 <= Compressor_14_3_F125_uid79_bh4_uid420_Out0(0);
   bh4_w18_10 <= Compressor_14_3_F125_uid79_bh4_uid420_Out0(1);
   bh4_w19_10 <= Compressor_14_3_F125_uid79_bh4_uid420_Out0(2);
   Compressor_14_3_F125_uid79_uid420: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid420_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid420_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid420_Out0_copy421);
   Compressor_14_3_F125_uid79_bh4_uid420_Out0 <= Compressor_14_3_F125_uid79_bh4_uid420_Out0_copy421; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid422_In0 <= "" & bh4_w19_9 & bh4_w19_8 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid422_In1 <= "" & bh4_w20_6;
   bh4_w19_11 <= Compressor_14_3_F125_uid79_bh4_uid422_Out0(0);
   bh4_w20_7 <= Compressor_14_3_F125_uid79_bh4_uid422_Out0(1);
   bh4_w21_8 <= Compressor_14_3_F125_uid79_bh4_uid422_Out0(2);
   Compressor_14_3_F125_uid79_uid422: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid422_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid422_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid422_Out0_copy423);
   Compressor_14_3_F125_uid79_bh4_uid422_Out0 <= Compressor_14_3_F125_uid79_bh4_uid422_Out0_copy423; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid424_In0 <= "" & bh4_w21_7 & bh4_w21_6 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid424_In1 <= "" & bh4_w22_6;
   bh4_w21_9 <= Compressor_14_3_F125_uid79_bh4_uid424_Out0(0);
   bh4_w22_7 <= Compressor_14_3_F125_uid79_bh4_uid424_Out0(1);
   bh4_w23_7 <= Compressor_14_3_F125_uid79_bh4_uid424_Out0(2);
   Compressor_14_3_F125_uid79_uid424: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid424_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid424_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid424_Out0_copy425);
   Compressor_14_3_F125_uid79_bh4_uid424_Out0 <= Compressor_14_3_F125_uid79_bh4_uid424_Out0_copy425; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid426_In0 <= "" & bh4_w23_6 & bh4_w23_5 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid426_In1 <= "" & bh4_w24_7;
   bh4_w23_8 <= Compressor_14_3_F125_uid79_bh4_uid426_Out0(0);
   bh4_w24_8 <= Compressor_14_3_F125_uid79_bh4_uid426_Out0(1);
   bh4_w25_6 <= Compressor_14_3_F125_uid79_bh4_uid426_Out0(2);
   Compressor_14_3_F125_uid79_uid426: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid426_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid426_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid426_Out0_copy427);
   Compressor_14_3_F125_uid79_bh4_uid426_Out0 <= Compressor_14_3_F125_uid79_bh4_uid426_Out0_copy427; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid428_In0 <= "" & bh4_w25_5 & bh4_w25_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid428_In1 <= "" & bh4_w26_8;
   bh4_w25_7 <= Compressor_14_3_F125_uid79_bh4_uid428_Out0(0);
   bh4_w26_9 <= Compressor_14_3_F125_uid79_bh4_uid428_Out0(1);
   bh4_w27_6 <= Compressor_14_3_F125_uid79_bh4_uid428_Out0(2);
   Compressor_14_3_F125_uid79_uid428: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid428_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid428_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid428_Out0_copy429);
   Compressor_14_3_F125_uid79_bh4_uid428_Out0 <= Compressor_14_3_F125_uid79_bh4_uid428_Out0_copy429; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid430_In0 <= "" & bh4_w28_9 & bh4_w28_8 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid430_In1 <= "" & bh4_w29_5;
   bh4_w28_10 <= Compressor_14_3_F125_uid79_bh4_uid430_Out0(0);
   bh4_w29_6 <= Compressor_14_3_F125_uid79_bh4_uid430_Out0(1);
   bh4_w30_10 <= Compressor_14_3_F125_uid79_bh4_uid430_Out0(2);
   Compressor_14_3_F125_uid79_uid430: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid430_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid430_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid430_Out0_copy431);
   Compressor_14_3_F125_uid79_bh4_uid430_Out0 <= Compressor_14_3_F125_uid79_bh4_uid430_Out0_copy431; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid432_In0 <= "" & bh4_w30_9 & bh4_w30_8 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid432_In1 <= "" & bh4_w31_5;
   bh4_w30_11 <= Compressor_14_3_F125_uid79_bh4_uid432_Out0(0);
   bh4_w31_6 <= Compressor_14_3_F125_uid79_bh4_uid432_Out0(1);
   bh4_w32_10 <= Compressor_14_3_F125_uid79_bh4_uid432_Out0(2);
   Compressor_14_3_F125_uid79_uid432: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid432_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid432_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid432_Out0_copy433);
   Compressor_14_3_F125_uid79_bh4_uid432_Out0 <= Compressor_14_3_F125_uid79_bh4_uid432_Out0_copy433; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid434_In0 <= "" & bh4_w32_9 & bh4_w32_8 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid434_In1 <= "" & bh4_w33_5;
   bh4_w32_11 <= Compressor_14_3_F125_uid79_bh4_uid434_Out0(0);
   bh4_w33_6 <= Compressor_14_3_F125_uid79_bh4_uid434_Out0(1);
   bh4_w34_10 <= Compressor_14_3_F125_uid79_bh4_uid434_Out0(2);
   Compressor_14_3_F125_uid79_uid434: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid434_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid434_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid434_Out0_copy435);
   Compressor_14_3_F125_uid79_bh4_uid434_Out0 <= Compressor_14_3_F125_uid79_bh4_uid434_Out0_copy435; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid436_In0 <= "" & bh4_w34_9 & bh4_w34_8 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid436_In1 <= "" & bh4_w35_5;
   bh4_w34_11 <= Compressor_14_3_F125_uid79_bh4_uid436_Out0(0);
   bh4_w35_6 <= Compressor_14_3_F125_uid79_bh4_uid436_Out0(1);
   bh4_w36_8 <= Compressor_14_3_F125_uid79_bh4_uid436_Out0(2);
   Compressor_14_3_F125_uid79_uid436: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid436_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid436_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid436_Out0_copy437);
   Compressor_14_3_F125_uid79_bh4_uid436_Out0 <= Compressor_14_3_F125_uid79_bh4_uid436_Out0_copy437; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid438_In0 <= "" & bh4_w36_7 & bh4_w36_6 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid438_In1 <= "" & bh4_w37_3;
   bh4_w36_9 <= Compressor_14_3_F125_uid79_bh4_uid438_Out0(0);
   bh4_w37_4 <= Compressor_14_3_F125_uid79_bh4_uid438_Out0(1);
   bh4_w38_6 <= Compressor_14_3_F125_uid79_bh4_uid438_Out0(2);
   Compressor_14_3_F125_uid79_uid438: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid438_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid438_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid438_Out0_copy439);
   Compressor_14_3_F125_uid79_bh4_uid438_Out0 <= Compressor_14_3_F125_uid79_bh4_uid438_Out0_copy439; -- output copy to hold a pipeline register if needed


   Compressor_14_3_F125_uid79_bh4_uid440_In0 <= "" & bh4_w38_5 & bh4_w38_4 & "0" & "0";
   Compressor_14_3_F125_uid79_bh4_uid440_In1 <= "" & bh4_w39_1;
   bh4_w38_7 <= Compressor_14_3_F125_uid79_bh4_uid440_Out0(0);
   bh4_w39_2 <= Compressor_14_3_F125_uid79_bh4_uid440_Out0(1);
   bh4_w40_1 <= Compressor_14_3_F125_uid79_bh4_uid440_Out0(2);
   Compressor_14_3_F125_uid79_uid440: Compressor_14_3_F125_uid79
      port map ( X0 => Compressor_14_3_F125_uid79_bh4_uid440_In0,
                 X1 => Compressor_14_3_F125_uid79_bh4_uid440_In1,
                 R => Compressor_14_3_F125_uid79_bh4_uid440_Out0_copy441);
   Compressor_14_3_F125_uid79_bh4_uid440_Out0 <= Compressor_14_3_F125_uid79_bh4_uid440_Out0_copy441; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh4_4 <= bh4_w4_60 & bh4_w3_59 & bh4_w2_54 & bh4_w1_45 & bh4_w0_34;

   bitheapFinalAdd_bh4_In0 <= "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & bh4_w40_1 & bh4_w39_2 & bh4_w38_7 & bh4_w37_4 & bh4_w36_9 & bh4_w35_6 & bh4_w34_11 & bh4_w33_6 & bh4_w32_11 & bh4_w31_6 & bh4_w30_11 & bh4_w29_6 & bh4_w28_10 & bh4_w27_6 & bh4_w26_9 & bh4_w25_7 & bh4_w24_8 & bh4_w23_8 & bh4_w22_7 & bh4_w21_9 & bh4_w20_7 & bh4_w19_11 & bh4_w18_10 & bh4_w17_15 & bh4_w16_15 & bh4_w15_23 & bh4_w14_24 & bh4_w13_30 & bh4_w12_33 & bh4_w11_36 & bh4_w10_39 & bh4_w9_43 & bh4_w8_46 & bh4_w7_53 & bh4_w6_56 & bh4_w5_59;
   bitheapFinalAdd_bh4_In1 <= "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & bh4_w40_0 & "0" & bh4_w38_6 & "0" & bh4_w36_8 & "0" & bh4_w34_10 & "0" & bh4_w32_10 & "0" & bh4_w30_10 & "0" & "0" & bh4_w27_5 & "0" & bh4_w25_6 & "0" & bh4_w23_7 & "0" & bh4_w21_8 & "0" & bh4_w19_10 & "0" & "0" & bh4_w16_14 & bh4_w15_22 & "0" & bh4_w13_29 & "0" & bh4_w11_35 & "0" & bh4_w9_42 & bh4_w8_44 & bh4_w7_52 & bh4_w6_55 & bh4_w5_58;
   bitheapFinalAdd_bh4_Cin <= '0';

   bitheapFinalAdd_bh4: IntAdder_64_F125_uid443
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh4_Cin,
                 X => bitheapFinalAdd_bh4_In0,
                 Y => bitheapFinalAdd_bh4_In1,
                 R => bitheapFinalAdd_bh4_Out);
   bitheapResult_bh4 <= bitheapFinalAdd_bh4_Out(62 downto 0) & tmp_bitheapResult_bh4_4;
   R <= bitheapResult_bh4(38 downto 5);
end architecture;
