-- Takes in one input (following AXI conventions), sending to four outputs at the same time.
library ieee;
use ieee.std_logic_1164.all;

entity axi_splitter_9 is
  generic (bit_width : natural);
  port ( clk        : in std_logic;
         rst      : in std_logic;

         in_ready_0 : out std_logic;
         in_valid_0 : in std_logic;
         in_data_0  : in std_logic_vector (bit_width-1 downto 0);

         out_ready_0 : in std_logic;
         out_valid_0 : out std_logic;
         out_data_0 : out std_logic_vector (bit_width-1 downto 0);

         out_ready_1 : in std_logic;
         out_valid_1 : out std_logic;
         out_data_1 : out std_logic_vector (bit_width-1 downto 0);

         out_ready_2 : in std_logic;
         out_valid_2 : out std_logic;
         out_data_2 : out std_logic_vector (bit_width-1 downto 0);

         out_ready_3 : in std_logic;
         out_valid_3 : out std_logic;
         out_data_3 : out std_logic_vector (bit_width-1 downto 0);

         out_ready_4 : in std_logic;
         out_valid_4 : out std_logic;
         out_data_4 : out std_logic_vector (bit_width-1 downto 0);

         out_ready_5 : in std_logic;
         out_valid_5 : out std_logic;
         out_data_5 : out std_logic_vector (bit_width-1 downto 0);

         out_ready_6 : in std_logic;
         out_valid_6 : out std_logic;
         out_data_6 : out std_logic_vector (bit_width-1 downto 0);

         out_ready_7 : in std_logic;
         out_valid_7 : out std_logic;
         out_data_7 : out std_logic_vector (bit_width-1 downto 0);

         out_ready_8 : in std_logic;
         out_valid_8 : out std_logic;
         out_data_8 : out std_logic_vector (bit_width-1 downto 0) );
end axi_splitter_9;

architecture Behavioral of axi_splitter_9 is
  signal temp_data_0   : std_logic_vector (bit_width-1 downto 0);
  signal is_in_ready_0 : std_logic := '1';
  signal is_stored_0   : std_logic := '0';
  signal is_sent       : std_logic := '0';

begin

  store_data : process(clk) -- store data when available in temporary storage
  begin
    if falling_edge(clk) then
      -- clear previous data (considered sent after 1 cycle where out valid and ready = 1)
      if (is_stored_0 = '1' AND (out_ready_0 = '1' AND out_ready_1 = '1' AND out_ready_2 = '1' AND out_ready_3 = '1' AND out_ready_4 = '1' AND out_ready_5 = '1' AND out_ready_6 = '1' AND out_ready_7 = '1' AND out_ready_8 = '1')) then
        is_stored_0 <= '0';
        is_in_ready_0 <= '1';
      else
        -- store data if input available and temp storage not used
        if (is_stored_0 = '0' AND
            in_valid_0 = '1' AND is_in_ready_0 = '1') then
          is_in_ready_0 <= '0';
          is_stored_0 <= '1';
          temp_data_0(bit_width-1 downto 0) <= in_data_0;
        end if;
      end if;
      -- for resetting component
      if (rst = '1') then
        is_stored_0 <= '0';
        is_in_ready_0 <= '1';
        is_sent <= '0';
      end if;
    end if;
  end process store_data;

  write_data : process(clk) -- write stored data to output ports
  begin
    if rising_edge(clk) then
      if (is_stored_0 = '1') then -- only write when both data ready to send
        out_data_0 <= temp_data_0(bit_width-1 downto 0);
        out_data_1 <= temp_data_0(bit_width-1 downto 0);
        out_data_2 <= temp_data_0(bit_width-1 downto 0);
        out_data_3 <= temp_data_0(bit_width-1 downto 0);
        out_data_4 <= temp_data_0(bit_width-1 downto 0);
        out_data_5 <= temp_data_0(bit_width-1 downto 0);
        out_data_6 <= temp_data_0(bit_width-1 downto 0);
        out_data_7 <= temp_data_0(bit_width-1 downto 0);
        out_data_8 <= temp_data_0(bit_width-1 downto 0);
      end if;
      in_ready_0 <= is_in_ready_0;
      out_valid_0 <= is_stored_0;
      out_valid_1 <= is_stored_0;
      out_valid_2 <= is_stored_0;
      out_valid_3 <= is_stored_0;
      out_valid_4 <= is_stored_0;
      out_valid_5 <= is_stored_0;
      out_valid_6 <= is_stored_0;
      out_valid_7 <= is_stored_0;
      out_valid_8 <= is_stored_0;
    end if;
  end process write_data;

end Behavioral;
